* File: acc_min_max.pex.sp
* Created: Tue Jan 16 15:28:05 2024
* Program "Calibre xRC"
* Version "v2016.4_15.11"
* 
.include "acc_min_max.pex.sp.pex"
.subckt acc_min_max_v3  VDD VSS ACC14 ACC12 ACC1 ACC11 ACC10 ACC9 ACC8 ACC7 ACC6
+ ACC5 ACC4 ACC3 ACC2 ACC0 ACC13 ACC15 MIN15 MIN14 MIN13 MIN12 MIN11 MIN10 MIN9
+ MIN8 MIN7 MIN6 MIN5 MIN4 MIN3 MIN2 MIN1 MIN0 CIN2 MAX15 MAX14 MAX13 MAX12
+ MAX11 MAX10 MAX9 MAX8 MAX7 MAX6 MAX5 MAX4 MAX3 MAX2 MAX1 MAX0 CIN1 Q CLEAR A15
+ A14 A13 A12 A11 A10 A9 A8 A7 A6 A5 A4 A3 A2 A1 A0 CLK
* 
* CLK	CLK
* A0	A0
* A1	A1
* A2	A2
* A3	A3
* A4	A4
* A5	A5
* A6	A6
* A7	A7
* A8	A8
* A9	A9
* A10	A10
* A11	A11
* A12	A12
* A13	A13
* A14	A14
* A15	A15
* CLEAR	CLEAR
* Q	Q
* CIN1	CIN1
* MAX0	MAX0
* MAX1	MAX1
* MAX2	MAX2
* MAX3	MAX3
* MAX4	MAX4
* MAX5	MAX5
* MAX6	MAX6
* MAX7	MAX7
* MAX8	MAX8
* MAX9	MAX9
* MAX10	MAX10
* MAX11	MAX11
* MAX12	MAX12
* MAX13	MAX13
* MAX14	MAX14
* MAX15	MAX15
* CIN2	CIN2
* MIN0	MIN0
* MIN1	MIN1
* MIN2	MIN2
* MIN3	MIN3
* MIN4	MIN4
* MIN5	MIN5
* MIN6	MIN6
* MIN7	MIN7
* MIN8	MIN8
* MIN9	MIN9
* MIN10	MIN10
* MIN11	MIN11
* MIN12	MIN12
* MIN13	MIN13
* MIN14	MIN14
* MIN15	MIN15
* ACC15	ACC15
* ACC13	ACC13
* ACC0	ACC0
* ACC2	ACC2
* ACC3	ACC3
* ACC4	ACC4
* ACC5	ACC5
* ACC6	ACC6
* ACC7	ACC7
* ACC8	ACC8
* ACC9	ACC9
* ACC10	ACC10
* ACC11	ACC11
* ACC1	ACC1
* ACC12	ACC12
* ACC14	ACC14
* VSS	VSS
* VDD	VDD
mXI10.XI0.XI0.MM2 N_XI10.XI0.NET0180_XI10.XI0.XI0.MM2_d
+ N_NET222_XI10.XI0.XI0.MM2_g N_VSS_XI10.XI0.XI0.MM2_s N_VSS_XI10.XI0.XI0.MM2_b
+ N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI10.XI0.XI1.MM2 N_XI10.XI0.NET35_XI10.XI0.XI1.MM2_d
+ N_XI10.XI0.NET0180_XI10.XI0.XI1.MM2_g N_VSS_XI10.XI0.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI25.MM2 N_NET206_XI25.MM2_d N_CLEAR_XI25.MM2_g N_VSS_XI25.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI24.MM2 N_NET202_XI24.MM2_d N_NET206_XI24.MM2_g N_VSS_XI24.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI23.XI11.MM2 N_NET696_XI23.XI11.MM2_d N_A15_XI23.XI11.MM2_g
+ N_VSS_XI23.XI11.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI22.XI11.MM2 N_NET662_XI22.XI11.MM2_d N_NET696_XI22.XI11.MM2_g
+ N_VSS_XI22.XI11.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI23.XI12.MM2 N_NET697_XI23.XI12.MM2_d N_A14_XI23.XI12.MM2_g
+ N_VSS_XI23.XI12.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI22.XI12.MM2 N_NET663_XI22.XI12.MM2_d N_NET697_XI22.XI12.MM2_g
+ N_VSS_XI22.XI12.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI23.XI10.MM2 N_NET698_XI23.XI10.MM2_d N_A13_XI23.XI10.MM2_g
+ N_VSS_XI23.XI10.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI22.XI10.MM2 N_NET664_XI22.XI10.MM2_d N_NET698_XI22.XI10.MM2_g
+ N_VSS_XI22.XI10.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI23.XI9.MM2 N_NET699_XI23.XI9.MM2_d N_A12_XI23.XI9.MM2_g N_VSS_XI23.XI9.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI22.XI9.MM2 N_NET665_XI22.XI9.MM2_d N_NET699_XI22.XI9.MM2_g
+ N_VSS_XI22.XI9.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI23.XI14.MM2 N_NET700_XI23.XI14.MM2_d N_A11_XI23.XI14.MM2_g
+ N_VSS_XI23.XI14.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI22.XI14.MM2 N_NET666_XI22.XI14.MM2_d N_NET700_XI22.XI14.MM2_g
+ N_VSS_XI22.XI14.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI23.XI13.MM2 N_NET701_XI23.XI13.MM2_d N_A10_XI23.XI13.MM2_g
+ N_VSS_XI23.XI13.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI22.XI13.MM2 N_NET667_XI22.XI13.MM2_d N_NET701_XI22.XI13.MM2_g
+ N_VSS_XI22.XI13.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI23.XI15.MM2 N_NET702_XI23.XI15.MM2_d N_A9_XI23.XI15.MM2_g
+ N_VSS_XI23.XI15.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI22.XI15.MM2 N_NET668_XI22.XI15.MM2_d N_NET702_XI22.XI15.MM2_g
+ N_VSS_XI22.XI15.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI23.XI6.MM2 N_NET703_XI23.XI6.MM2_d N_A8_XI23.XI6.MM2_g N_VSS_XI23.XI6.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI22.XI6.MM2 N_NET669_XI22.XI6.MM2_d N_NET703_XI22.XI6.MM2_g
+ N_VSS_XI22.XI6.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI23.XI5.MM2 N_NET704_XI23.XI5.MM2_d N_A7_XI23.XI5.MM2_g N_VSS_XI23.XI5.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI22.XI5.MM2 N_NET670_XI22.XI5.MM2_d N_NET704_XI22.XI5.MM2_g
+ N_VSS_XI22.XI5.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI23.XI7.MM2 N_NET705_XI23.XI7.MM2_d N_A6_XI23.XI7.MM2_g N_VSS_XI23.XI7.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI22.XI7.MM2 N_NET671_XI22.XI7.MM2_d N_NET705_XI22.XI7.MM2_g
+ N_VSS_XI22.XI7.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI23.XI8.MM2 N_NET706_XI23.XI8.MM2_d N_A5_XI23.XI8.MM2_g N_VSS_XI23.XI8.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI22.XI8.MM2 N_NET672_XI22.XI8.MM2_d N_NET706_XI22.XI8.MM2_g
+ N_VSS_XI22.XI8.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI23.XI3.MM2 N_NET707_XI23.XI3.MM2_d N_A4_XI23.XI3.MM2_g N_VSS_XI23.XI3.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI22.XI3.MM2 N_NET673_XI22.XI3.MM2_d N_NET707_XI22.XI3.MM2_g
+ N_VSS_XI22.XI3.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI23.XI4.MM2 N_NET708_XI23.XI4.MM2_d N_A3_XI23.XI4.MM2_g N_VSS_XI23.XI4.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI22.XI4.MM2 N_NET674_XI22.XI4.MM2_d N_NET708_XI22.XI4.MM2_g
+ N_VSS_XI22.XI4.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI23.XI2.MM2 N_NET709_XI23.XI2.MM2_d N_A2_XI23.XI2.MM2_g N_VSS_XI23.XI2.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI22.XI2.MM2 N_NET675_XI22.XI2.MM2_d N_NET709_XI22.XI2.MM2_g
+ N_VSS_XI22.XI2.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI23.XI1.MM2 N_NET710_XI23.XI1.MM2_d N_A1_XI23.XI1.MM2_g N_VSS_XI23.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI22.XI1.MM2 N_NET676_XI22.XI1.MM2_d N_NET710_XI22.XI1.MM2_g
+ N_VSS_XI22.XI1.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI23.XI0.MM2 N_NET711_XI23.XI0.MM2_d N_A0_XI23.XI0.MM2_g N_VSS_XI23.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI22.XI0.MM2 N_NET677_XI22.XI0.MM2_d N_NET711_XI22.XI0.MM2_g
+ N_VSS_XI22.XI0.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI10.XI0.MM26 N_XI10.XI0.CLKB_XI10.XI0.MM26_d N_XI10.XI0.NET35_XI10.XI0.MM26_g
+ N_VSS_XI10.XI0.MM26_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI17.XI0.MM2 N_XI17.NET0180_XI17.XI0.MM2_d N_NET222_XI17.XI0.MM2_g
+ N_VSS_XI17.XI0.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI17.XI1.MM2 N_XI17.NET35_XI17.XI1.MM2_d N_XI17.NET0180_XI17.XI1.MM2_g
+ N_VSS_XI17.XI1.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI17.MM26 N_XI17.CLKB_XI17.MM26_d N_XI17.NET35_XI17.MM26_g N_VSS_XI17.MM26_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI17.MM19 N_XI17.NET27_XI17.MM19_d N_NET202_XI17.MM19_g N_VSS_XI17.MM19_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI17.MM18 N_XI17.NET31_XI17.MM18_d N_XI17.NET27_XI17.MM18_g N_VSS_XI17.MM18_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI17.MM28 N_XI17.NET31_XI17.MM28_d N_XI17.CLKB_XI17.MM28_g
+ N_XI17.NET58_XI17.MM28_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI17.MM6 N_XI17.NET15_XI17.MM6_d N_XI17.NET58_XI17.MM6_g N_VSS_XI17.MM6_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI17.MM0 N_XI17.NET54_XI17.MM0_d N_XI17.NET15_XI17.MM0_g N_VSS_XI17.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI17.MM36 N_XI17.NET58_XI17.MM36_d N_XI17.NET35_XI17.MM36_g
+ N_XI17.NET54_XI17.MM36_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI17.MM38 N_XI17.NET15_XI17.MM38_d N_XI17.NET35_XI17.MM38_g
+ N_XI17.NET14_XI17.MM38_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI17.MM15 N_Q_XI17.MM15_d N_XI17.NET14_XI17.MM15_g N_VSS_XI17.MM15_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI17.MM16 N_NET198_XI17.MM16_d N_Q_XI17.MM16_g N_VSS_XI17.MM16_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI17.MM40 N_XI17.NET14_XI17.MM40_d N_XI17.CLKB_XI17.MM40_g N_NET198_XI17.MM40_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI0.MM19 N_XI10.XI0.NET27_XI10.XI0.MM19_d N_NET677_XI10.XI0.MM19_g
+ N_VSS_XI10.XI0.MM19_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI10.XI0.MM18 N_XI10.XI0.NET31_XI10.XI0.MM18_d N_XI10.XI0.NET27_XI10.XI0.MM18_g
+ N_VSS_XI10.XI0.MM18_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI10.XI30.XI0.MM2 N_XI10.XI30.NET0180_XI10.XI30.XI0.MM2_d
+ N_NET222_XI10.XI30.XI0.MM2_g N_VSS_XI10.XI30.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI29.XI0.MM2 N_XI10.XI29.NET0180_XI10.XI29.XI0.MM2_d
+ N_NET222_XI10.XI29.XI0.MM2_g N_VSS_XI10.XI29.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI31.XI0.MM2 N_XI10.XI31.NET0180_XI10.XI31.XI0.MM2_d
+ N_NET222_XI10.XI31.XI0.MM2_g N_VSS_XI10.XI31.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI28.XI0.MM2 N_XI10.XI28.NET0180_XI10.XI28.XI0.MM2_d
+ N_NET222_XI10.XI28.XI0.MM2_g N_VSS_XI10.XI28.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI25.XI0.MM2 N_XI10.XI25.NET0180_XI10.XI25.XI0.MM2_d
+ N_NET222_XI10.XI25.XI0.MM2_g N_VSS_XI10.XI25.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI26.XI0.MM2 N_XI10.XI26.NET0180_XI10.XI26.XI0.MM2_d
+ N_NET222_XI10.XI26.XI0.MM2_g N_VSS_XI10.XI26.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI24.XI0.MM2 N_XI10.XI24.NET0180_XI10.XI24.XI0.MM2_d
+ N_NET222_XI10.XI24.XI0.MM2_g N_VSS_XI10.XI24.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI27.XI0.MM2 N_XI10.XI27.NET0180_XI10.XI27.XI0.MM2_d
+ N_NET222_XI10.XI27.XI0.MM2_g N_VSS_XI10.XI27.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI22.XI0.MM2 N_XI10.XI22.NET0180_XI10.XI22.XI0.MM2_d
+ N_NET222_XI10.XI22.XI0.MM2_g N_VSS_XI10.XI22.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI21.XI0.MM2 N_XI10.XI21.NET0180_XI10.XI21.XI0.MM2_d
+ N_NET222_XI10.XI21.XI0.MM2_g N_VSS_XI10.XI21.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI23.XI0.MM2 N_XI10.XI23.NET0180_XI10.XI23.XI0.MM2_d
+ N_NET222_XI10.XI23.XI0.MM2_g N_VSS_XI10.XI23.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI19.XI0.MM2 N_XI10.XI19.NET0180_XI10.XI19.XI0.MM2_d
+ N_NET222_XI10.XI19.XI0.MM2_g N_VSS_XI10.XI19.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI20.XI0.MM2 N_XI10.XI20.NET0180_XI10.XI20.XI0.MM2_d
+ N_NET222_XI10.XI20.XI0.MM2_g N_VSS_XI10.XI20.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI18.XI0.MM2 N_XI10.XI18.NET0180_XI10.XI18.XI0.MM2_d
+ N_NET222_XI10.XI18.XI0.MM2_g N_VSS_XI10.XI18.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI17.XI0.MM2 N_XI10.XI17.NET0180_XI10.XI17.XI0.MM2_d
+ N_NET222_XI10.XI17.XI0.MM2_g N_VSS_XI10.XI17.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI0.MM28 N_XI10.XI0.NET31_XI10.XI0.MM28_d N_XI10.XI0.CLKB_XI10.XI0.MM28_g
+ N_XI10.XI0.NET58_XI10.XI0.MM28_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI10.XI30.XI1.MM2 N_XI10.XI30.NET35_XI10.XI30.XI1.MM2_d
+ N_XI10.XI30.NET0180_XI10.XI30.XI1.MM2_g N_VSS_XI10.XI30.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI29.XI1.MM2 N_XI10.XI29.NET35_XI10.XI29.XI1.MM2_d
+ N_XI10.XI29.NET0180_XI10.XI29.XI1.MM2_g N_VSS_XI10.XI29.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI31.XI1.MM2 N_XI10.XI31.NET35_XI10.XI31.XI1.MM2_d
+ N_XI10.XI31.NET0180_XI10.XI31.XI1.MM2_g N_VSS_XI10.XI31.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI28.XI1.MM2 N_XI10.XI28.NET35_XI10.XI28.XI1.MM2_d
+ N_XI10.XI28.NET0180_XI10.XI28.XI1.MM2_g N_VSS_XI10.XI28.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI25.XI1.MM2 N_XI10.XI25.NET35_XI10.XI25.XI1.MM2_d
+ N_XI10.XI25.NET0180_XI10.XI25.XI1.MM2_g N_VSS_XI10.XI25.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI26.XI1.MM2 N_XI10.XI26.NET35_XI10.XI26.XI1.MM2_d
+ N_XI10.XI26.NET0180_XI10.XI26.XI1.MM2_g N_VSS_XI10.XI26.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI24.XI1.MM2 N_XI10.XI24.NET35_XI10.XI24.XI1.MM2_d
+ N_XI10.XI24.NET0180_XI10.XI24.XI1.MM2_g N_VSS_XI10.XI24.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI27.XI1.MM2 N_XI10.XI27.NET35_XI10.XI27.XI1.MM2_d
+ N_XI10.XI27.NET0180_XI10.XI27.XI1.MM2_g N_VSS_XI10.XI27.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI22.XI1.MM2 N_XI10.XI22.NET35_XI10.XI22.XI1.MM2_d
+ N_XI10.XI22.NET0180_XI10.XI22.XI1.MM2_g N_VSS_XI10.XI22.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI21.XI1.MM2 N_XI10.XI21.NET35_XI10.XI21.XI1.MM2_d
+ N_XI10.XI21.NET0180_XI10.XI21.XI1.MM2_g N_VSS_XI10.XI21.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI23.XI1.MM2 N_XI10.XI23.NET35_XI10.XI23.XI1.MM2_d
+ N_XI10.XI23.NET0180_XI10.XI23.XI1.MM2_g N_VSS_XI10.XI23.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI19.XI1.MM2 N_XI10.XI19.NET35_XI10.XI19.XI1.MM2_d
+ N_XI10.XI19.NET0180_XI10.XI19.XI1.MM2_g N_VSS_XI10.XI19.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI20.XI1.MM2 N_XI10.XI20.NET35_XI10.XI20.XI1.MM2_d
+ N_XI10.XI20.NET0180_XI10.XI20.XI1.MM2_g N_VSS_XI10.XI20.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI18.XI1.MM2 N_XI10.XI18.NET35_XI10.XI18.XI1.MM2_d
+ N_XI10.XI18.NET0180_XI10.XI18.XI1.MM2_g N_VSS_XI10.XI18.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI17.XI1.MM2 N_XI10.XI17.NET35_XI10.XI17.XI1.MM2_d
+ N_XI10.XI17.NET0180_XI10.XI17.XI1.MM2_g N_VSS_XI10.XI17.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI0.MM6 N_XI10.XI0.NET15_XI10.XI0.MM6_d N_XI10.XI0.NET58_XI10.XI0.MM6_g
+ N_VSS_XI10.XI0.MM6_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI10.XI30.MM26 N_XI10.XI30.CLKB_XI10.XI30.MM26_d
+ N_XI10.XI30.NET35_XI10.XI30.MM26_g N_VSS_XI10.XI30.MM26_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI29.MM26 N_XI10.XI29.CLKB_XI10.XI29.MM26_d
+ N_XI10.XI29.NET35_XI10.XI29.MM26_g N_VSS_XI10.XI29.MM26_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI31.MM26 N_XI10.XI31.CLKB_XI10.XI31.MM26_d
+ N_XI10.XI31.NET35_XI10.XI31.MM26_g N_VSS_XI10.XI31.MM26_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI28.MM26 N_XI10.XI28.CLKB_XI10.XI28.MM26_d
+ N_XI10.XI28.NET35_XI10.XI28.MM26_g N_VSS_XI10.XI28.MM26_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI25.MM26 N_XI10.XI25.CLKB_XI10.XI25.MM26_d
+ N_XI10.XI25.NET35_XI10.XI25.MM26_g N_VSS_XI10.XI25.MM26_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI26.MM26 N_XI10.XI26.CLKB_XI10.XI26.MM26_d
+ N_XI10.XI26.NET35_XI10.XI26.MM26_g N_VSS_XI10.XI26.MM26_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI24.MM26 N_XI10.XI24.CLKB_XI10.XI24.MM26_d
+ N_XI10.XI24.NET35_XI10.XI24.MM26_g N_VSS_XI10.XI24.MM26_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI27.MM26 N_XI10.XI27.CLKB_XI10.XI27.MM26_d
+ N_XI10.XI27.NET35_XI10.XI27.MM26_g N_VSS_XI10.XI27.MM26_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI22.MM26 N_XI10.XI22.CLKB_XI10.XI22.MM26_d
+ N_XI10.XI22.NET35_XI10.XI22.MM26_g N_VSS_XI10.XI22.MM26_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI21.MM26 N_XI10.XI21.CLKB_XI10.XI21.MM26_d
+ N_XI10.XI21.NET35_XI10.XI21.MM26_g N_VSS_XI10.XI21.MM26_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI23.MM26 N_XI10.XI23.CLKB_XI10.XI23.MM26_d
+ N_XI10.XI23.NET35_XI10.XI23.MM26_g N_VSS_XI10.XI23.MM26_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI19.MM26 N_XI10.XI19.CLKB_XI10.XI19.MM26_d
+ N_XI10.XI19.NET35_XI10.XI19.MM26_g N_VSS_XI10.XI19.MM26_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI20.MM26 N_XI10.XI20.CLKB_XI10.XI20.MM26_d
+ N_XI10.XI20.NET35_XI10.XI20.MM26_g N_VSS_XI10.XI20.MM26_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI18.MM26 N_XI10.XI18.CLKB_XI10.XI18.MM26_d
+ N_XI10.XI18.NET35_XI10.XI18.MM26_g N_VSS_XI10.XI18.MM26_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI17.MM26 N_XI10.XI17.CLKB_XI10.XI17.MM26_d
+ N_XI10.XI17.NET35_XI10.XI17.MM26_g N_VSS_XI10.XI17.MM26_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI0.MM0 N_XI10.XI0.NET54_XI10.XI0.MM0_d N_XI10.XI0.NET15_XI10.XI0.MM0_g
+ N_VSS_XI10.XI0.MM0_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI10.XI30.MM19 N_XI10.XI30.NET27_XI10.XI30.MM19_d N_NET662_XI10.XI30.MM19_g
+ N_VSS_XI10.XI30.MM19_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI10.XI29.MM19 N_XI10.XI29.NET27_XI10.XI29.MM19_d N_NET663_XI10.XI29.MM19_g
+ N_VSS_XI10.XI29.MM19_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI10.XI31.MM19 N_XI10.XI31.NET27_XI10.XI31.MM19_d N_NET664_XI10.XI31.MM19_g
+ N_VSS_XI10.XI31.MM19_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI10.XI28.MM19 N_XI10.XI28.NET27_XI10.XI28.MM19_d N_NET665_XI10.XI28.MM19_g
+ N_VSS_XI10.XI28.MM19_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI10.XI25.MM19 N_XI10.XI25.NET27_XI10.XI25.MM19_d N_NET666_XI10.XI25.MM19_g
+ N_VSS_XI10.XI25.MM19_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI10.XI26.MM19 N_XI10.XI26.NET27_XI10.XI26.MM19_d N_NET667_XI10.XI26.MM19_g
+ N_VSS_XI10.XI26.MM19_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI10.XI24.MM19 N_XI10.XI24.NET27_XI10.XI24.MM19_d N_NET668_XI10.XI24.MM19_g
+ N_VSS_XI10.XI24.MM19_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI10.XI27.MM19 N_XI10.XI27.NET27_XI10.XI27.MM19_d N_NET669_XI10.XI27.MM19_g
+ N_VSS_XI10.XI27.MM19_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI10.XI22.MM19 N_XI10.XI22.NET27_XI10.XI22.MM19_d N_NET670_XI10.XI22.MM19_g
+ N_VSS_XI10.XI22.MM19_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI10.XI21.MM19 N_XI10.XI21.NET27_XI10.XI21.MM19_d N_NET671_XI10.XI21.MM19_g
+ N_VSS_XI10.XI21.MM19_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI10.XI23.MM19 N_XI10.XI23.NET27_XI10.XI23.MM19_d N_NET672_XI10.XI23.MM19_g
+ N_VSS_XI10.XI23.MM19_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI10.XI19.MM19 N_XI10.XI19.NET27_XI10.XI19.MM19_d N_NET673_XI10.XI19.MM19_g
+ N_VSS_XI10.XI19.MM19_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI10.XI20.MM19 N_XI10.XI20.NET27_XI10.XI20.MM19_d N_NET674_XI10.XI20.MM19_g
+ N_VSS_XI10.XI20.MM19_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI10.XI18.MM19 N_XI10.XI18.NET27_XI10.XI18.MM19_d N_NET675_XI10.XI18.MM19_g
+ N_VSS_XI10.XI18.MM19_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI10.XI17.MM19 N_XI10.XI17.NET27_XI10.XI17.MM19_d N_NET676_XI10.XI17.MM19_g
+ N_VSS_XI10.XI17.MM19_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI10.XI0.MM36 N_XI10.XI0.NET58_XI10.XI0.MM36_d N_XI10.XI0.NET35_XI10.XI0.MM36_g
+ N_XI10.XI0.NET54_XI10.XI0.MM36_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI10.XI30.MM18 N_XI10.XI30.NET31_XI10.XI30.MM18_d
+ N_XI10.XI30.NET27_XI10.XI30.MM18_g N_VSS_XI10.XI30.MM18_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI29.MM18 N_XI10.XI29.NET31_XI10.XI29.MM18_d
+ N_XI10.XI29.NET27_XI10.XI29.MM18_g N_VSS_XI10.XI29.MM18_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI31.MM18 N_XI10.XI31.NET31_XI10.XI31.MM18_d
+ N_XI10.XI31.NET27_XI10.XI31.MM18_g N_VSS_XI10.XI31.MM18_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI28.MM18 N_XI10.XI28.NET31_XI10.XI28.MM18_d
+ N_XI10.XI28.NET27_XI10.XI28.MM18_g N_VSS_XI10.XI28.MM18_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI25.MM18 N_XI10.XI25.NET31_XI10.XI25.MM18_d
+ N_XI10.XI25.NET27_XI10.XI25.MM18_g N_VSS_XI10.XI25.MM18_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI26.MM18 N_XI10.XI26.NET31_XI10.XI26.MM18_d
+ N_XI10.XI26.NET27_XI10.XI26.MM18_g N_VSS_XI10.XI26.MM18_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI24.MM18 N_XI10.XI24.NET31_XI10.XI24.MM18_d
+ N_XI10.XI24.NET27_XI10.XI24.MM18_g N_VSS_XI10.XI24.MM18_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI27.MM18 N_XI10.XI27.NET31_XI10.XI27.MM18_d
+ N_XI10.XI27.NET27_XI10.XI27.MM18_g N_VSS_XI10.XI27.MM18_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI22.MM18 N_XI10.XI22.NET31_XI10.XI22.MM18_d
+ N_XI10.XI22.NET27_XI10.XI22.MM18_g N_VSS_XI10.XI22.MM18_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI21.MM18 N_XI10.XI21.NET31_XI10.XI21.MM18_d
+ N_XI10.XI21.NET27_XI10.XI21.MM18_g N_VSS_XI10.XI21.MM18_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI23.MM18 N_XI10.XI23.NET31_XI10.XI23.MM18_d
+ N_XI10.XI23.NET27_XI10.XI23.MM18_g N_VSS_XI10.XI23.MM18_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI19.MM18 N_XI10.XI19.NET31_XI10.XI19.MM18_d
+ N_XI10.XI19.NET27_XI10.XI19.MM18_g N_VSS_XI10.XI19.MM18_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI20.MM18 N_XI10.XI20.NET31_XI10.XI20.MM18_d
+ N_XI10.XI20.NET27_XI10.XI20.MM18_g N_VSS_XI10.XI20.MM18_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI18.MM18 N_XI10.XI18.NET31_XI10.XI18.MM18_d
+ N_XI10.XI18.NET27_XI10.XI18.MM18_g N_VSS_XI10.XI18.MM18_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI17.MM18 N_XI10.XI17.NET31_XI10.XI17.MM18_d
+ N_XI10.XI17.NET27_XI10.XI17.MM18_g N_VSS_XI10.XI17.MM18_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI0.MM38 N_XI10.XI0.NET15_XI10.XI0.MM38_d N_XI10.XI0.NET35_XI10.XI0.MM38_g
+ N_XI10.XI0.NET14_XI10.XI0.MM38_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI10.XI30.MM28 N_XI10.XI30.NET31_XI10.XI30.MM28_d
+ N_XI10.XI30.CLKB_XI10.XI30.MM28_g N_XI10.XI30.NET58_XI10.XI30.MM28_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI29.MM28 N_XI10.XI29.NET31_XI10.XI29.MM28_d
+ N_XI10.XI29.CLKB_XI10.XI29.MM28_g N_XI10.XI29.NET58_XI10.XI29.MM28_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI31.MM28 N_XI10.XI31.NET31_XI10.XI31.MM28_d
+ N_XI10.XI31.CLKB_XI10.XI31.MM28_g N_XI10.XI31.NET58_XI10.XI31.MM28_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI28.MM28 N_XI10.XI28.NET31_XI10.XI28.MM28_d
+ N_XI10.XI28.CLKB_XI10.XI28.MM28_g N_XI10.XI28.NET58_XI10.XI28.MM28_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI25.MM28 N_XI10.XI25.NET31_XI10.XI25.MM28_d
+ N_XI10.XI25.CLKB_XI10.XI25.MM28_g N_XI10.XI25.NET58_XI10.XI25.MM28_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI26.MM28 N_XI10.XI26.NET31_XI10.XI26.MM28_d
+ N_XI10.XI26.CLKB_XI10.XI26.MM28_g N_XI10.XI26.NET58_XI10.XI26.MM28_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI24.MM28 N_XI10.XI24.NET31_XI10.XI24.MM28_d
+ N_XI10.XI24.CLKB_XI10.XI24.MM28_g N_XI10.XI24.NET58_XI10.XI24.MM28_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI27.MM28 N_XI10.XI27.NET31_XI10.XI27.MM28_d
+ N_XI10.XI27.CLKB_XI10.XI27.MM28_g N_XI10.XI27.NET58_XI10.XI27.MM28_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI22.MM28 N_XI10.XI22.NET31_XI10.XI22.MM28_d
+ N_XI10.XI22.CLKB_XI10.XI22.MM28_g N_XI10.XI22.NET58_XI10.XI22.MM28_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI21.MM28 N_XI10.XI21.NET31_XI10.XI21.MM28_d
+ N_XI10.XI21.CLKB_XI10.XI21.MM28_g N_XI10.XI21.NET58_XI10.XI21.MM28_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI23.MM28 N_XI10.XI23.NET31_XI10.XI23.MM28_d
+ N_XI10.XI23.CLKB_XI10.XI23.MM28_g N_XI10.XI23.NET58_XI10.XI23.MM28_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI19.MM28 N_XI10.XI19.NET31_XI10.XI19.MM28_d
+ N_XI10.XI19.CLKB_XI10.XI19.MM28_g N_XI10.XI19.NET58_XI10.XI19.MM28_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI20.MM28 N_XI10.XI20.NET31_XI10.XI20.MM28_d
+ N_XI10.XI20.CLKB_XI10.XI20.MM28_g N_XI10.XI20.NET58_XI10.XI20.MM28_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI18.MM28 N_XI10.XI18.NET31_XI10.XI18.MM28_d
+ N_XI10.XI18.CLKB_XI10.XI18.MM28_g N_XI10.XI18.NET58_XI10.XI18.MM28_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI17.MM28 N_XI10.XI17.NET31_XI10.XI17.MM28_d
+ N_XI10.XI17.CLKB_XI10.XI17.MM28_g N_XI10.XI17.NET58_XI10.XI17.MM28_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI0.MM15 N_NET256_XI10.XI0.MM15_d N_XI10.XI0.NET14_XI10.XI0.MM15_g
+ N_VSS_XI10.XI0.MM15_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI10.XI30.MM6 N_XI10.XI30.NET15_XI10.XI30.MM6_d
+ N_XI10.XI30.NET58_XI10.XI30.MM6_g N_VSS_XI10.XI30.MM6_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI29.MM6 N_XI10.XI29.NET15_XI10.XI29.MM6_d
+ N_XI10.XI29.NET58_XI10.XI29.MM6_g N_VSS_XI10.XI29.MM6_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI31.MM6 N_XI10.XI31.NET15_XI10.XI31.MM6_d
+ N_XI10.XI31.NET58_XI10.XI31.MM6_g N_VSS_XI10.XI31.MM6_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI28.MM6 N_XI10.XI28.NET15_XI10.XI28.MM6_d
+ N_XI10.XI28.NET58_XI10.XI28.MM6_g N_VSS_XI10.XI28.MM6_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI25.MM6 N_XI10.XI25.NET15_XI10.XI25.MM6_d
+ N_XI10.XI25.NET58_XI10.XI25.MM6_g N_VSS_XI10.XI25.MM6_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI26.MM6 N_XI10.XI26.NET15_XI10.XI26.MM6_d
+ N_XI10.XI26.NET58_XI10.XI26.MM6_g N_VSS_XI10.XI26.MM6_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI24.MM6 N_XI10.XI24.NET15_XI10.XI24.MM6_d
+ N_XI10.XI24.NET58_XI10.XI24.MM6_g N_VSS_XI10.XI24.MM6_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI27.MM6 N_XI10.XI27.NET15_XI10.XI27.MM6_d
+ N_XI10.XI27.NET58_XI10.XI27.MM6_g N_VSS_XI10.XI27.MM6_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI22.MM6 N_XI10.XI22.NET15_XI10.XI22.MM6_d
+ N_XI10.XI22.NET58_XI10.XI22.MM6_g N_VSS_XI10.XI22.MM6_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI21.MM6 N_XI10.XI21.NET15_XI10.XI21.MM6_d
+ N_XI10.XI21.NET58_XI10.XI21.MM6_g N_VSS_XI10.XI21.MM6_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI23.MM6 N_XI10.XI23.NET15_XI10.XI23.MM6_d
+ N_XI10.XI23.NET58_XI10.XI23.MM6_g N_VSS_XI10.XI23.MM6_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI19.MM6 N_XI10.XI19.NET15_XI10.XI19.MM6_d
+ N_XI10.XI19.NET58_XI10.XI19.MM6_g N_VSS_XI10.XI19.MM6_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI20.MM6 N_XI10.XI20.NET15_XI10.XI20.MM6_d
+ N_XI10.XI20.NET58_XI10.XI20.MM6_g N_VSS_XI10.XI20.MM6_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI18.MM6 N_XI10.XI18.NET15_XI10.XI18.MM6_d
+ N_XI10.XI18.NET58_XI10.XI18.MM6_g N_VSS_XI10.XI18.MM6_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI17.MM6 N_XI10.XI17.NET15_XI10.XI17.MM6_d
+ N_XI10.XI17.NET58_XI10.XI17.MM6_g N_VSS_XI10.XI17.MM6_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI0.MM16 N_XI10.BAR_Q1_XI10.XI0.MM16_d N_NET256_XI10.XI0.MM16_g
+ N_VSS_XI10.XI0.MM16_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI10.XI30.MM0 N_XI10.XI30.NET54_XI10.XI30.MM0_d
+ N_XI10.XI30.NET15_XI10.XI30.MM0_g N_VSS_XI10.XI30.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI29.MM0 N_XI10.XI29.NET54_XI10.XI29.MM0_d
+ N_XI10.XI29.NET15_XI10.XI29.MM0_g N_VSS_XI10.XI29.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI31.MM0 N_XI10.XI31.NET54_XI10.XI31.MM0_d
+ N_XI10.XI31.NET15_XI10.XI31.MM0_g N_VSS_XI10.XI31.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI28.MM0 N_XI10.XI28.NET54_XI10.XI28.MM0_d
+ N_XI10.XI28.NET15_XI10.XI28.MM0_g N_VSS_XI10.XI28.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI25.MM0 N_XI10.XI25.NET54_XI10.XI25.MM0_d
+ N_XI10.XI25.NET15_XI10.XI25.MM0_g N_VSS_XI10.XI25.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI26.MM0 N_XI10.XI26.NET54_XI10.XI26.MM0_d
+ N_XI10.XI26.NET15_XI10.XI26.MM0_g N_VSS_XI10.XI26.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI24.MM0 N_XI10.XI24.NET54_XI10.XI24.MM0_d
+ N_XI10.XI24.NET15_XI10.XI24.MM0_g N_VSS_XI10.XI24.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI27.MM0 N_XI10.XI27.NET54_XI10.XI27.MM0_d
+ N_XI10.XI27.NET15_XI10.XI27.MM0_g N_VSS_XI10.XI27.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI22.MM0 N_XI10.XI22.NET54_XI10.XI22.MM0_d
+ N_XI10.XI22.NET15_XI10.XI22.MM0_g N_VSS_XI10.XI22.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI21.MM0 N_XI10.XI21.NET54_XI10.XI21.MM0_d
+ N_XI10.XI21.NET15_XI10.XI21.MM0_g N_VSS_XI10.XI21.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI23.MM0 N_XI10.XI23.NET54_XI10.XI23.MM0_d
+ N_XI10.XI23.NET15_XI10.XI23.MM0_g N_VSS_XI10.XI23.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI19.MM0 N_XI10.XI19.NET54_XI10.XI19.MM0_d
+ N_XI10.XI19.NET15_XI10.XI19.MM0_g N_VSS_XI10.XI19.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI20.MM0 N_XI10.XI20.NET54_XI10.XI20.MM0_d
+ N_XI10.XI20.NET15_XI10.XI20.MM0_g N_VSS_XI10.XI20.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI18.MM0 N_XI10.XI18.NET54_XI10.XI18.MM0_d
+ N_XI10.XI18.NET15_XI10.XI18.MM0_g N_VSS_XI10.XI18.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI17.MM0 N_XI10.XI17.NET54_XI10.XI17.MM0_d
+ N_XI10.XI17.NET15_XI10.XI17.MM0_g N_VSS_XI10.XI17.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI0.MM40 N_XI10.XI0.NET14_XI10.XI0.MM40_d N_XI10.XI0.CLKB_XI10.XI0.MM40_g
+ N_XI10.BAR_Q1_XI10.XI0.MM40_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI10.XI30.MM36 N_XI10.XI30.NET58_XI10.XI30.MM36_d
+ N_XI10.XI30.NET35_XI10.XI30.MM36_g N_XI10.XI30.NET54_XI10.XI30.MM36_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI29.MM36 N_XI10.XI29.NET58_XI10.XI29.MM36_d
+ N_XI10.XI29.NET35_XI10.XI29.MM36_g N_XI10.XI29.NET54_XI10.XI29.MM36_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI31.MM36 N_XI10.XI31.NET58_XI10.XI31.MM36_d
+ N_XI10.XI31.NET35_XI10.XI31.MM36_g N_XI10.XI31.NET54_XI10.XI31.MM36_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI28.MM36 N_XI10.XI28.NET58_XI10.XI28.MM36_d
+ N_XI10.XI28.NET35_XI10.XI28.MM36_g N_XI10.XI28.NET54_XI10.XI28.MM36_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI25.MM36 N_XI10.XI25.NET58_XI10.XI25.MM36_d
+ N_XI10.XI25.NET35_XI10.XI25.MM36_g N_XI10.XI25.NET54_XI10.XI25.MM36_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI26.MM36 N_XI10.XI26.NET58_XI10.XI26.MM36_d
+ N_XI10.XI26.NET35_XI10.XI26.MM36_g N_XI10.XI26.NET54_XI10.XI26.MM36_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI24.MM36 N_XI10.XI24.NET58_XI10.XI24.MM36_d
+ N_XI10.XI24.NET35_XI10.XI24.MM36_g N_XI10.XI24.NET54_XI10.XI24.MM36_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI27.MM36 N_XI10.XI27.NET58_XI10.XI27.MM36_d
+ N_XI10.XI27.NET35_XI10.XI27.MM36_g N_XI10.XI27.NET54_XI10.XI27.MM36_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI22.MM36 N_XI10.XI22.NET58_XI10.XI22.MM36_d
+ N_XI10.XI22.NET35_XI10.XI22.MM36_g N_XI10.XI22.NET54_XI10.XI22.MM36_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI21.MM36 N_XI10.XI21.NET58_XI10.XI21.MM36_d
+ N_XI10.XI21.NET35_XI10.XI21.MM36_g N_XI10.XI21.NET54_XI10.XI21.MM36_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI23.MM36 N_XI10.XI23.NET58_XI10.XI23.MM36_d
+ N_XI10.XI23.NET35_XI10.XI23.MM36_g N_XI10.XI23.NET54_XI10.XI23.MM36_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI19.MM36 N_XI10.XI19.NET58_XI10.XI19.MM36_d
+ N_XI10.XI19.NET35_XI10.XI19.MM36_g N_XI10.XI19.NET54_XI10.XI19.MM36_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI20.MM36 N_XI10.XI20.NET58_XI10.XI20.MM36_d
+ N_XI10.XI20.NET35_XI10.XI20.MM36_g N_XI10.XI20.NET54_XI10.XI20.MM36_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI18.MM36 N_XI10.XI18.NET58_XI10.XI18.MM36_d
+ N_XI10.XI18.NET35_XI10.XI18.MM36_g N_XI10.XI18.NET54_XI10.XI18.MM36_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI17.MM36 N_XI10.XI17.NET58_XI10.XI17.MM36_d
+ N_XI10.XI17.NET35_XI10.XI17.MM36_g N_XI10.XI17.NET54_XI10.XI17.MM36_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI30.MM38 N_XI10.XI30.NET15_XI10.XI30.MM38_d
+ N_XI10.XI30.NET35_XI10.XI30.MM38_g N_XI10.XI30.NET14_XI10.XI30.MM38_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI29.MM38 N_XI10.XI29.NET15_XI10.XI29.MM38_d
+ N_XI10.XI29.NET35_XI10.XI29.MM38_g N_XI10.XI29.NET14_XI10.XI29.MM38_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI31.MM38 N_XI10.XI31.NET15_XI10.XI31.MM38_d
+ N_XI10.XI31.NET35_XI10.XI31.MM38_g N_XI10.XI31.NET14_XI10.XI31.MM38_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI28.MM38 N_XI10.XI28.NET15_XI10.XI28.MM38_d
+ N_XI10.XI28.NET35_XI10.XI28.MM38_g N_XI10.XI28.NET14_XI10.XI28.MM38_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI25.MM38 N_XI10.XI25.NET15_XI10.XI25.MM38_d
+ N_XI10.XI25.NET35_XI10.XI25.MM38_g N_XI10.XI25.NET14_XI10.XI25.MM38_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI26.MM38 N_XI10.XI26.NET15_XI10.XI26.MM38_d
+ N_XI10.XI26.NET35_XI10.XI26.MM38_g N_XI10.XI26.NET14_XI10.XI26.MM38_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI24.MM38 N_XI10.XI24.NET15_XI10.XI24.MM38_d
+ N_XI10.XI24.NET35_XI10.XI24.MM38_g N_XI10.XI24.NET14_XI10.XI24.MM38_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI27.MM38 N_XI10.XI27.NET15_XI10.XI27.MM38_d
+ N_XI10.XI27.NET35_XI10.XI27.MM38_g N_XI10.XI27.NET14_XI10.XI27.MM38_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI22.MM38 N_XI10.XI22.NET15_XI10.XI22.MM38_d
+ N_XI10.XI22.NET35_XI10.XI22.MM38_g N_XI10.XI22.NET14_XI10.XI22.MM38_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI21.MM38 N_XI10.XI21.NET15_XI10.XI21.MM38_d
+ N_XI10.XI21.NET35_XI10.XI21.MM38_g N_XI10.XI21.NET14_XI10.XI21.MM38_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI23.MM38 N_XI10.XI23.NET15_XI10.XI23.MM38_d
+ N_XI10.XI23.NET35_XI10.XI23.MM38_g N_XI10.XI23.NET14_XI10.XI23.MM38_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI19.MM38 N_XI10.XI19.NET15_XI10.XI19.MM38_d
+ N_XI10.XI19.NET35_XI10.XI19.MM38_g N_XI10.XI19.NET14_XI10.XI19.MM38_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI20.MM38 N_XI10.XI20.NET15_XI10.XI20.MM38_d
+ N_XI10.XI20.NET35_XI10.XI20.MM38_g N_XI10.XI20.NET14_XI10.XI20.MM38_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI18.MM38 N_XI10.XI18.NET15_XI10.XI18.MM38_d
+ N_XI10.XI18.NET35_XI10.XI18.MM38_g N_XI10.XI18.NET14_XI10.XI18.MM38_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI17.MM38 N_XI10.XI17.NET15_XI10.XI17.MM38_d
+ N_XI10.XI17.NET35_XI10.XI17.MM38_g N_XI10.XI17.NET14_XI10.XI17.MM38_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI9.XI97.XI4.MM2 N_XI9.XI97.NET39_XI9.XI97.XI4.MM2_d N_CIN1_XI9.XI97.XI4.MM2_g
+ N_VSS_XI9.XI97.XI4.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI10.XI30.MM15 N_NET241_XI10.XI30.MM15_d N_XI10.XI30.NET14_XI10.XI30.MM15_g
+ N_VSS_XI10.XI30.MM15_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI10.XI29.MM15 N_NET242_XI10.XI29.MM15_d N_XI10.XI29.NET14_XI10.XI29.MM15_g
+ N_VSS_XI10.XI29.MM15_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI10.XI31.MM15 N_NET243_XI10.XI31.MM15_d N_XI10.XI31.NET14_XI10.XI31.MM15_g
+ N_VSS_XI10.XI31.MM15_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI10.XI28.MM15 N_NET244_XI10.XI28.MM15_d N_XI10.XI28.NET14_XI10.XI28.MM15_g
+ N_VSS_XI10.XI28.MM15_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI10.XI25.MM15 N_NET245_XI10.XI25.MM15_d N_XI10.XI25.NET14_XI10.XI25.MM15_g
+ N_VSS_XI10.XI25.MM15_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI10.XI26.MM15 N_NET246_XI10.XI26.MM15_d N_XI10.XI26.NET14_XI10.XI26.MM15_g
+ N_VSS_XI10.XI26.MM15_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI10.XI24.MM15 N_NET247_XI10.XI24.MM15_d N_XI10.XI24.NET14_XI10.XI24.MM15_g
+ N_VSS_XI10.XI24.MM15_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI10.XI27.MM15 N_NET248_XI10.XI27.MM15_d N_XI10.XI27.NET14_XI10.XI27.MM15_g
+ N_VSS_XI10.XI27.MM15_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI10.XI22.MM15 N_NET249_XI10.XI22.MM15_d N_XI10.XI22.NET14_XI10.XI22.MM15_g
+ N_VSS_XI10.XI22.MM15_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI10.XI21.MM15 N_NET250_XI10.XI21.MM15_d N_XI10.XI21.NET14_XI10.XI21.MM15_g
+ N_VSS_XI10.XI21.MM15_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI10.XI23.MM15 N_NET251_XI10.XI23.MM15_d N_XI10.XI23.NET14_XI10.XI23.MM15_g
+ N_VSS_XI10.XI23.MM15_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI10.XI19.MM15 N_NET252_XI10.XI19.MM15_d N_XI10.XI19.NET14_XI10.XI19.MM15_g
+ N_VSS_XI10.XI19.MM15_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI10.XI20.MM15 N_NET253_XI10.XI20.MM15_d N_XI10.XI20.NET14_XI10.XI20.MM15_g
+ N_VSS_XI10.XI20.MM15_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI10.XI18.MM15 N_NET254_XI10.XI18.MM15_d N_XI10.XI18.NET14_XI10.XI18.MM15_g
+ N_VSS_XI10.XI18.MM15_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI10.XI17.MM15 N_NET255_XI10.XI17.MM15_d N_XI10.XI17.NET14_XI10.XI17.MM15_g
+ N_VSS_XI10.XI17.MM15_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI9.XI97.MM7 N_XI9.XI97.NET10_XI9.XI97.MM7_d N_XI9.XI97.NET39_XI9.XI97.MM7_g
+ N_VSS_XI9.XI97.MM7_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.2375e-13 AS=3.225e-13 PD=8.95e-07 PS=1.79e-06
mXI9.XI97.MM2 N_NET192_XI9.XI97.MM2_d N_XI9.XI97.NET43_XI9.XI97.MM2_g
+ N_XI9.XI97.NET10_XI9.XI97.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=4.75e-13 AS=2.2375e-13 PD=1.9e-06 PS=8.95e-07
mXI10.XI30.MM16 N_XI10.BAR_Q16_XI10.XI30.MM16_d N_NET241_XI10.XI30.MM16_g
+ N_VSS_XI10.XI30.MM16_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI10.XI29.MM16 N_XI10.BAR_Q15_XI10.XI29.MM16_d N_NET242_XI10.XI29.MM16_g
+ N_VSS_XI10.XI29.MM16_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI10.XI31.MM16 N_XI10.BAR_Q14_XI10.XI31.MM16_d N_NET243_XI10.XI31.MM16_g
+ N_VSS_XI10.XI31.MM16_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI10.XI28.MM16 N_XI10.BAR_Q13_XI10.XI28.MM16_d N_NET244_XI10.XI28.MM16_g
+ N_VSS_XI10.XI28.MM16_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI10.XI25.MM16 N_XI10.BAR_Q12_XI10.XI25.MM16_d N_NET245_XI10.XI25.MM16_g
+ N_VSS_XI10.XI25.MM16_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI10.XI26.MM16 N_XI10.BAR_Q11_XI10.XI26.MM16_d N_NET246_XI10.XI26.MM16_g
+ N_VSS_XI10.XI26.MM16_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI10.XI24.MM16 N_XI10.BAR_Q10_XI10.XI24.MM16_d N_NET247_XI10.XI24.MM16_g
+ N_VSS_XI10.XI24.MM16_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI10.XI27.MM16 N_XI10.BAR_Q9_XI10.XI27.MM16_d N_NET248_XI10.XI27.MM16_g
+ N_VSS_XI10.XI27.MM16_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI10.XI22.MM16 N_XI10.BAR_Q8_XI10.XI22.MM16_d N_NET249_XI10.XI22.MM16_g
+ N_VSS_XI10.XI22.MM16_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI10.XI21.MM16 N_XI10.BAR_Q7_XI10.XI21.MM16_d N_NET250_XI10.XI21.MM16_g
+ N_VSS_XI10.XI21.MM16_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI10.XI23.MM16 N_XI10.BAR_Q6_XI10.XI23.MM16_d N_NET251_XI10.XI23.MM16_g
+ N_VSS_XI10.XI23.MM16_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI10.XI19.MM16 N_XI10.BAR_Q5_XI10.XI19.MM16_d N_NET252_XI10.XI19.MM16_g
+ N_VSS_XI10.XI19.MM16_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI10.XI20.MM16 N_XI10.BAR_Q4_XI10.XI20.MM16_d N_NET253_XI10.XI20.MM16_g
+ N_VSS_XI10.XI20.MM16_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI10.XI18.MM16 N_XI10.BAR_Q3_XI10.XI18.MM16_d N_NET254_XI10.XI18.MM16_g
+ N_VSS_XI10.XI18.MM16_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI10.XI17.MM16 N_XI10.BAR_Q2_XI10.XI17.MM16_d N_NET255_XI10.XI17.MM16_g
+ N_VSS_XI10.XI17.MM16_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI9.XI97.MM0 N_NET192_XI9.XI97.MM0_d N_XI9.P1_XI9.XI97.MM0_g
+ N_XI9.XI97.NET6_XI9.XI97.MM0_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=4.75e-13 AS=1.8125e-13 PD=1.9e-06 PS=7.25e-07
mXI10.XI30.MM40 N_XI10.XI30.NET14_XI10.XI30.MM40_d
+ N_XI10.XI30.CLKB_XI10.XI30.MM40_g N_XI10.BAR_Q16_XI10.XI30.MM40_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI29.MM40 N_XI10.XI29.NET14_XI10.XI29.MM40_d
+ N_XI10.XI29.CLKB_XI10.XI29.MM40_g N_XI10.BAR_Q15_XI10.XI29.MM40_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI31.MM40 N_XI10.XI31.NET14_XI10.XI31.MM40_d
+ N_XI10.XI31.CLKB_XI10.XI31.MM40_g N_XI10.BAR_Q14_XI10.XI31.MM40_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI28.MM40 N_XI10.XI28.NET14_XI10.XI28.MM40_d
+ N_XI10.XI28.CLKB_XI10.XI28.MM40_g N_XI10.BAR_Q13_XI10.XI28.MM40_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI25.MM40 N_XI10.XI25.NET14_XI10.XI25.MM40_d
+ N_XI10.XI25.CLKB_XI10.XI25.MM40_g N_XI10.BAR_Q12_XI10.XI25.MM40_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI26.MM40 N_XI10.XI26.NET14_XI10.XI26.MM40_d
+ N_XI10.XI26.CLKB_XI10.XI26.MM40_g N_XI10.BAR_Q11_XI10.XI26.MM40_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI24.MM40 N_XI10.XI24.NET14_XI10.XI24.MM40_d
+ N_XI10.XI24.CLKB_XI10.XI24.MM40_g N_XI10.BAR_Q10_XI10.XI24.MM40_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI27.MM40 N_XI10.XI27.NET14_XI10.XI27.MM40_d
+ N_XI10.XI27.CLKB_XI10.XI27.MM40_g N_XI10.BAR_Q9_XI10.XI27.MM40_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI22.MM40 N_XI10.XI22.NET14_XI10.XI22.MM40_d
+ N_XI10.XI22.CLKB_XI10.XI22.MM40_g N_XI10.BAR_Q8_XI10.XI22.MM40_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI21.MM40 N_XI10.XI21.NET14_XI10.XI21.MM40_d
+ N_XI10.XI21.CLKB_XI10.XI21.MM40_g N_XI10.BAR_Q7_XI10.XI21.MM40_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI23.MM40 N_XI10.XI23.NET14_XI10.XI23.MM40_d
+ N_XI10.XI23.CLKB_XI10.XI23.MM40_g N_XI10.BAR_Q6_XI10.XI23.MM40_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI19.MM40 N_XI10.XI19.NET14_XI10.XI19.MM40_d
+ N_XI10.XI19.CLKB_XI10.XI19.MM40_g N_XI10.BAR_Q5_XI10.XI19.MM40_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI20.MM40 N_XI10.XI20.NET14_XI10.XI20.MM40_d
+ N_XI10.XI20.CLKB_XI10.XI20.MM40_g N_XI10.BAR_Q4_XI10.XI20.MM40_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI18.MM40 N_XI10.XI18.NET14_XI10.XI18.MM40_d
+ N_XI10.XI18.CLKB_XI10.XI18.MM40_g N_XI10.BAR_Q3_XI10.XI18.MM40_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI10.XI17.MM40 N_XI10.XI17.NET14_XI10.XI17.MM40_d
+ N_XI10.XI17.CLKB_XI10.XI17.MM40_g N_XI10.BAR_Q2_XI10.XI17.MM40_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI9.XI97.MM6 N_XI9.XI97.NET6_XI9.XI97.MM6_d N_CIN1_XI9.XI97.MM6_g
+ N_VSS_XI9.XI97.MM6_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=1.8125e-13 AS=2.575e-13 PD=7.25e-07 PS=1.53e-06
mXI9.XI97.XI9.MM2 N_XI9.XI97.NET43_XI9.XI97.XI9.MM2_d
+ N_XI9.P1_XI9.XI97.XI9.MM2_g N_VSS_XI9.XI97.XI9.MM2_s N_VSS_XI10.XI0.XI0.MM2_b
+ N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9.XI153.XI1.MM0 N_XI9.XI153.XI1.NET036_XI9.XI153.XI1.MM0_d
+ N_NET242_XI9.XI153.XI1.MM0_g N_VSS_XI9.XI153.XI1.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.85e-13 AS=2.45e-13
+ PD=7.4e-07 PS=1.48e-06
mXI9.XI154.XI1.MM0 N_XI9.XI154.XI1.NET036_XI9.XI154.XI1.MM0_d
+ N_NET243_XI9.XI154.XI1.MM0_g N_VSS_XI9.XI154.XI1.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.85e-13 AS=2.45e-13
+ PD=7.4e-07 PS=1.48e-06
mXI9.XI157.XI1.MM0 N_XI9.XI157.XI1.NET036_XI9.XI157.XI1.MM0_d
+ N_NET244_XI9.XI157.XI1.MM0_g N_VSS_XI9.XI157.XI1.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.85e-13 AS=2.45e-13
+ PD=7.4e-07 PS=1.48e-06
mXI9.XI156.XI1.MM0 N_XI9.XI156.XI1.NET036_XI9.XI156.XI1.MM0_d
+ N_NET245_XI9.XI156.XI1.MM0_g N_VSS_XI9.XI156.XI1.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.85e-13 AS=2.45e-13
+ PD=7.4e-07 PS=1.48e-06
mXI9.XI155.XI1.MM0 N_XI9.XI155.XI1.NET036_XI9.XI155.XI1.MM0_d
+ N_NET246_XI9.XI155.XI1.MM0_g N_VSS_XI9.XI155.XI1.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.85e-13 AS=2.45e-13
+ PD=7.4e-07 PS=1.48e-06
mXI9.XI133.XI1.MM0 N_XI9.XI133.XI1.NET036_XI9.XI133.XI1.MM0_d
+ N_NET247_XI9.XI133.XI1.MM0_g N_VSS_XI9.XI133.XI1.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.85e-13 AS=2.45e-13
+ PD=7.4e-07 PS=1.48e-06
mXI9.XI132.XI1.MM0 N_XI9.XI132.XI1.NET036_XI9.XI132.XI1.MM0_d
+ N_NET248_XI9.XI132.XI1.MM0_g N_VSS_XI9.XI132.XI1.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.85e-13 AS=2.45e-13
+ PD=7.4e-07 PS=1.48e-06
mXI9.XI131.XI1.MM0 N_XI9.XI131.XI1.NET036_XI9.XI131.XI1.MM0_d
+ N_NET249_XI9.XI131.XI1.MM0_g N_VSS_XI9.XI131.XI1.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.85e-13 AS=2.45e-13
+ PD=7.4e-07 PS=1.48e-06
mXI9.XI111.XI1.MM0 N_XI9.XI111.XI1.NET036_XI9.XI111.XI1.MM0_d
+ N_NET250_XI9.XI111.XI1.MM0_g N_VSS_XI9.XI111.XI1.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.85e-13 AS=2.45e-13
+ PD=7.4e-07 PS=1.48e-06
mXI9.XI110.XI1.MM0 N_XI9.XI110.XI1.NET036_XI9.XI110.XI1.MM0_d
+ N_NET251_XI9.XI110.XI1.MM0_g N_VSS_XI9.XI110.XI1.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.85e-13 AS=2.45e-13
+ PD=7.4e-07 PS=1.48e-06
mXI9.XI103.XI1.MM0 N_XI9.XI103.XI1.NET036_XI9.XI103.XI1.MM0_d
+ N_NET252_XI9.XI103.XI1.MM0_g N_VSS_XI9.XI103.XI1.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.85e-13 AS=2.45e-13
+ PD=7.4e-07 PS=1.48e-06
mXI9.XI102.XI1.MM0 N_XI9.XI102.XI1.NET036_XI9.XI102.XI1.MM0_d
+ N_NET253_XI9.XI102.XI1.MM0_g N_VSS_XI9.XI102.XI1.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.85e-13 AS=2.45e-13
+ PD=7.4e-07 PS=1.48e-06
mXI9.XI88.XI1.MM0 N_XI9.XI88.XI1.NET036_XI9.XI88.XI1.MM0_d
+ N_NET254_XI9.XI88.XI1.MM0_g N_VSS_XI9.XI88.XI1.MM0_s N_VSS_XI10.XI0.XI0.MM2_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.85e-13 AS=2.45e-13 PD=7.4e-07 PS=1.48e-06
mXI9.XI82.XI1.MM0 N_XI9.XI82.XI1.NET036_XI9.XI82.XI1.MM0_d
+ N_NET255_XI9.XI82.XI1.MM0_g N_VSS_XI9.XI82.XI1.MM0_s N_VSS_XI10.XI0.XI0.MM2_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.85e-13 AS=2.45e-13 PD=7.4e-07 PS=1.48e-06
mXI9.XI10.XI1.MM0 N_XI9.XI10.XI1.NET036_XI9.XI10.XI1.MM0_d
+ N_NET256_XI9.XI10.XI1.MM0_g N_VSS_XI9.XI10.XI1.MM0_s N_VSS_XI10.XI0.XI0.MM2_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.85e-13 AS=2.45e-13 PD=7.4e-07 PS=1.48e-06
mXI9.XI153.XI1.MM2 N_XI9.XI153.NET6_XI9.XI153.XI1.MM2_d
+ N_ACC14_XI9.XI153.XI1.MM2_g N_XI9.XI153.XI1.NET036_XI9.XI153.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=1.85e-13
+ PD=1.52e-06 PS=7.4e-07
mXI9.XI154.XI1.MM2 N_XI9.XI154.NET6_XI9.XI154.XI1.MM2_d
+ N_ACC13_XI9.XI154.XI1.MM2_g N_XI9.XI154.XI1.NET036_XI9.XI154.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=1.85e-13
+ PD=1.52e-06 PS=7.4e-07
mXI9.XI157.XI1.MM2 N_XI9.XI157.NET6_XI9.XI157.XI1.MM2_d
+ N_ACC12_XI9.XI157.XI1.MM2_g N_XI9.XI157.XI1.NET036_XI9.XI157.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=1.85e-13
+ PD=1.52e-06 PS=7.4e-07
mXI9.XI156.XI1.MM2 N_XI9.XI156.NET6_XI9.XI156.XI1.MM2_d
+ N_ACC11_XI9.XI156.XI1.MM2_g N_XI9.XI156.XI1.NET036_XI9.XI156.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=1.85e-13
+ PD=1.52e-06 PS=7.4e-07
mXI9.XI155.XI1.MM2 N_XI9.XI155.NET6_XI9.XI155.XI1.MM2_d
+ N_ACC10_XI9.XI155.XI1.MM2_g N_XI9.XI155.XI1.NET036_XI9.XI155.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=1.85e-13
+ PD=1.52e-06 PS=7.4e-07
mXI9.XI133.XI1.MM2 N_XI9.XI133.NET6_XI9.XI133.XI1.MM2_d
+ N_ACC9_XI9.XI133.XI1.MM2_g N_XI9.XI133.XI1.NET036_XI9.XI133.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=1.85e-13
+ PD=1.52e-06 PS=7.4e-07
mXI9.XI132.XI1.MM2 N_XI9.XI132.NET6_XI9.XI132.XI1.MM2_d
+ N_ACC8_XI9.XI132.XI1.MM2_g N_XI9.XI132.XI1.NET036_XI9.XI132.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=1.85e-13
+ PD=1.52e-06 PS=7.4e-07
mXI9.XI131.XI1.MM2 N_XI9.XI131.NET6_XI9.XI131.XI1.MM2_d
+ N_ACC7_XI9.XI131.XI1.MM2_g N_XI9.XI131.XI1.NET036_XI9.XI131.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=1.85e-13
+ PD=1.52e-06 PS=7.4e-07
mXI9.XI111.XI1.MM2 N_XI9.XI111.NET6_XI9.XI111.XI1.MM2_d
+ N_ACC6_XI9.XI111.XI1.MM2_g N_XI9.XI111.XI1.NET036_XI9.XI111.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=1.85e-13
+ PD=1.52e-06 PS=7.4e-07
mXI9.XI110.XI1.MM2 N_XI9.XI110.NET6_XI9.XI110.XI1.MM2_d
+ N_ACC5_XI9.XI110.XI1.MM2_g N_XI9.XI110.XI1.NET036_XI9.XI110.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=1.85e-13
+ PD=1.52e-06 PS=7.4e-07
mXI9.XI103.XI1.MM2 N_XI9.XI103.NET6_XI9.XI103.XI1.MM2_d
+ N_ACC4_XI9.XI103.XI1.MM2_g N_XI9.XI103.XI1.NET036_XI9.XI103.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=1.85e-13
+ PD=1.52e-06 PS=7.4e-07
mXI9.XI102.XI1.MM2 N_XI9.XI102.NET6_XI9.XI102.XI1.MM2_d
+ N_ACC3_XI9.XI102.XI1.MM2_g N_XI9.XI102.XI1.NET036_XI9.XI102.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=1.85e-13
+ PD=1.52e-06 PS=7.4e-07
mXI9.XI88.XI1.MM2 N_XI9.XI88.NET6_XI9.XI88.XI1.MM2_d N_ACC2_XI9.XI88.XI1.MM2_g
+ N_XI9.XI88.XI1.NET036_XI9.XI88.XI1.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18
+ L=1.8e-07 W=5e-07 AD=2.55e-13 AS=1.85e-13 PD=1.52e-06 PS=7.4e-07
mXI9.XI82.XI1.MM2 N_XI9.XI82.NET6_XI9.XI82.XI1.MM2_d N_ACC1_XI9.XI82.XI1.MM2_g
+ N_XI9.XI82.XI1.NET036_XI9.XI82.XI1.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18
+ L=1.8e-07 W=5e-07 AD=2.55e-13 AS=1.85e-13 PD=1.52e-06 PS=7.4e-07
mXI9.XI10.XI1.MM2 N_XI9.XI10.NET6_XI9.XI10.XI1.MM2_d N_ACC0_XI9.XI10.XI1.MM2_g
+ N_XI9.XI10.XI1.NET036_XI9.XI10.XI1.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18
+ L=1.8e-07 W=5e-07 AD=2.55e-13 AS=1.85e-13 PD=1.52e-06 PS=7.4e-07
mXI9.XI134.XI4.MM2 N_XI9.XI134.NET39_XI9.XI134.XI4.MM2_d
+ N_NET241_XI9.XI134.XI4.MM2_g N_VSS_XI9.XI134.XI4.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI9.XI153.XI0.MM2 N_XI9.G15_XI9.XI153.XI0.MM2_d
+ N_XI9.XI153.NET6_XI9.XI153.XI0.MM2_g N_VSS_XI9.XI153.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI9.XI154.XI0.MM2 N_XI9.G14_XI9.XI154.XI0.MM2_d
+ N_XI9.XI154.NET6_XI9.XI154.XI0.MM2_g N_VSS_XI9.XI154.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI9.XI157.XI0.MM2 N_XI9.G13_XI9.XI157.XI0.MM2_d
+ N_XI9.XI157.NET6_XI9.XI157.XI0.MM2_g N_VSS_XI9.XI157.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI9.XI156.XI0.MM2 N_XI9.G12_XI9.XI156.XI0.MM2_d
+ N_XI9.XI156.NET6_XI9.XI156.XI0.MM2_g N_VSS_XI9.XI156.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI9.XI155.XI0.MM2 N_XI9.G11_XI9.XI155.XI0.MM2_d
+ N_XI9.XI155.NET6_XI9.XI155.XI0.MM2_g N_VSS_XI9.XI155.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI9.XI133.XI0.MM2 N_XI9.G10_XI9.XI133.XI0.MM2_d
+ N_XI9.XI133.NET6_XI9.XI133.XI0.MM2_g N_VSS_XI9.XI133.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI9.XI132.XI0.MM2 N_XI9.G9_XI9.XI132.XI0.MM2_d
+ N_XI9.XI132.NET6_XI9.XI132.XI0.MM2_g N_VSS_XI9.XI132.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI9.XI131.XI0.MM2 N_XI9.G8_XI9.XI131.XI0.MM2_d
+ N_XI9.XI131.NET6_XI9.XI131.XI0.MM2_g N_VSS_XI9.XI131.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI9.XI111.XI0.MM2 N_XI9.G7_XI9.XI111.XI0.MM2_d
+ N_XI9.XI111.NET6_XI9.XI111.XI0.MM2_g N_VSS_XI9.XI111.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI9.XI110.XI0.MM2 N_XI9.G6_XI9.XI110.XI0.MM2_d
+ N_XI9.XI110.NET6_XI9.XI110.XI0.MM2_g N_VSS_XI9.XI110.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI9.XI103.XI0.MM2 N_XI9.G5_XI9.XI103.XI0.MM2_d
+ N_XI9.XI103.NET6_XI9.XI103.XI0.MM2_g N_VSS_XI9.XI103.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI9.XI102.XI0.MM2 N_XI9.G4_XI9.XI102.XI0.MM2_d
+ N_XI9.XI102.NET6_XI9.XI102.XI0.MM2_g N_VSS_XI9.XI102.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI9.XI88.XI0.MM2 N_XI9.G3_XI9.XI88.XI0.MM2_d N_XI9.XI88.NET6_XI9.XI88.XI0.MM2_g
+ N_VSS_XI9.XI88.XI0.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9.XI82.XI0.MM2 N_XI9.G2_XI9.XI82.XI0.MM2_d N_XI9.XI82.NET6_XI9.XI82.XI0.MM2_g
+ N_VSS_XI9.XI82.XI0.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9.XI10.XI0.MM2 N_XI9.G1_XI9.XI10.XI0.MM2_d N_XI9.XI10.NET6_XI9.XI10.XI0.MM2_g
+ N_VSS_XI9.XI10.XI0.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9.XI134.MM7 N_XI9.XI134.NET10_XI9.XI134.MM7_d
+ N_XI9.XI134.NET39_XI9.XI134.MM7_g N_VSS_XI9.XI134.MM7_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.2375e-13 AS=3.225e-13
+ PD=8.95e-07 PS=1.79e-06
mXI9.XI134.MM2 N_XI9.P16_XI9.XI134.MM2_d N_XI9.XI134.NET43_XI9.XI134.MM2_g
+ N_XI9.XI134.NET10_XI9.XI134.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=4.75e-13 AS=2.2375e-13 PD=1.9e-06 PS=8.95e-07
mXI9.XI137.XI4.MM2 N_XI9.XI137.NET39_XI9.XI137.XI4.MM2_d
+ N_NET242_XI9.XI137.XI4.MM2_g N_VSS_XI9.XI137.XI4.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI9.XI140.XI4.MM2 N_XI9.XI140.NET39_XI9.XI140.XI4.MM2_d
+ N_NET243_XI9.XI140.XI4.MM2_g N_VSS_XI9.XI140.XI4.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI9.XI149.XI4.MM2 N_XI9.XI149.NET39_XI9.XI149.XI4.MM2_d
+ N_NET244_XI9.XI149.XI4.MM2_g N_VSS_XI9.XI149.XI4.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI9.XI146.XI4.MM2 N_XI9.XI146.NET39_XI9.XI146.XI4.MM2_d
+ N_NET245_XI9.XI146.XI4.MM2_g N_VSS_XI9.XI146.XI4.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI9.XI143.XI4.MM2 N_XI9.XI143.NET39_XI9.XI143.XI4.MM2_d
+ N_NET246_XI9.XI143.XI4.MM2_g N_VSS_XI9.XI143.XI4.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI9.XI128.XI4.MM2 N_XI9.XI128.NET39_XI9.XI128.XI4.MM2_d
+ N_NET247_XI9.XI128.XI4.MM2_g N_VSS_XI9.XI128.XI4.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI9.XI125.XI4.MM2 N_XI9.XI125.NET39_XI9.XI125.XI4.MM2_d
+ N_NET248_XI9.XI125.XI4.MM2_g N_VSS_XI9.XI125.XI4.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI9.XI122.XI4.MM2 N_XI9.XI122.NET39_XI9.XI122.XI4.MM2_d
+ N_NET249_XI9.XI122.XI4.MM2_g N_VSS_XI9.XI122.XI4.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI9.XI114.XI4.MM2 N_XI9.XI114.NET39_XI9.XI114.XI4.MM2_d
+ N_NET250_XI9.XI114.XI4.MM2_g N_VSS_XI9.XI114.XI4.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI9.XI109.XI4.MM2 N_XI9.XI109.NET39_XI9.XI109.XI4.MM2_d
+ N_NET251_XI9.XI109.XI4.MM2_g N_VSS_XI9.XI109.XI4.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI9.XI106.XI4.MM2 N_XI9.XI106.NET39_XI9.XI106.XI4.MM2_d
+ N_NET252_XI9.XI106.XI4.MM2_g N_VSS_XI9.XI106.XI4.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI9.XI101.XI4.MM2 N_XI9.XI101.NET39_XI9.XI101.XI4.MM2_d
+ N_NET253_XI9.XI101.XI4.MM2_g N_VSS_XI9.XI101.XI4.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI9.XI86.XI4.MM2 N_XI9.XI86.NET39_XI9.XI86.XI4.MM2_d
+ N_NET254_XI9.XI86.XI4.MM2_g N_VSS_XI9.XI86.XI4.MM2_s N_VSS_XI10.XI0.XI0.MM2_b
+ N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9.XI80.XI4.MM2 N_XI9.XI80.NET39_XI9.XI80.XI4.MM2_d
+ N_NET255_XI9.XI80.XI4.MM2_g N_VSS_XI9.XI80.XI4.MM2_s N_VSS_XI10.XI0.XI0.MM2_b
+ N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9.XI26.XI4.MM2 N_XI9.XI26.NET39_XI9.XI26.XI4.MM2_d
+ N_NET256_XI9.XI26.XI4.MM2_g N_VSS_XI9.XI26.XI4.MM2_s N_VSS_XI10.XI0.XI0.MM2_b
+ N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9.XI134.MM0 N_XI9.P16_XI9.XI134.MM0_d N_ACC15_XI9.XI134.MM0_g
+ N_XI9.XI134.NET6_XI9.XI134.MM0_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=4.75e-13 AS=1.8125e-13 PD=1.9e-06 PS=7.25e-07
mXI9.XI137.MM7 N_XI9.XI137.NET10_XI9.XI137.MM7_d
+ N_XI9.XI137.NET39_XI9.XI137.MM7_g N_VSS_XI9.XI137.MM7_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.2375e-13 AS=3.225e-13
+ PD=8.95e-07 PS=1.79e-06
mXI9.XI140.MM7 N_XI9.XI140.NET10_XI9.XI140.MM7_d
+ N_XI9.XI140.NET39_XI9.XI140.MM7_g N_VSS_XI9.XI140.MM7_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.2375e-13 AS=3.225e-13
+ PD=8.95e-07 PS=1.79e-06
mXI9.XI149.MM7 N_XI9.XI149.NET10_XI9.XI149.MM7_d
+ N_XI9.XI149.NET39_XI9.XI149.MM7_g N_VSS_XI9.XI149.MM7_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.2375e-13 AS=3.225e-13
+ PD=8.95e-07 PS=1.79e-06
mXI9.XI146.MM7 N_XI9.XI146.NET10_XI9.XI146.MM7_d
+ N_XI9.XI146.NET39_XI9.XI146.MM7_g N_VSS_XI9.XI146.MM7_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.2375e-13 AS=3.225e-13
+ PD=8.95e-07 PS=1.79e-06
mXI9.XI143.MM7 N_XI9.XI143.NET10_XI9.XI143.MM7_d
+ N_XI9.XI143.NET39_XI9.XI143.MM7_g N_VSS_XI9.XI143.MM7_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.2375e-13 AS=3.225e-13
+ PD=8.95e-07 PS=1.79e-06
mXI9.XI128.MM7 N_XI9.XI128.NET10_XI9.XI128.MM7_d
+ N_XI9.XI128.NET39_XI9.XI128.MM7_g N_VSS_XI9.XI128.MM7_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.2375e-13 AS=3.225e-13
+ PD=8.95e-07 PS=1.79e-06
mXI9.XI125.MM7 N_XI9.XI125.NET10_XI9.XI125.MM7_d
+ N_XI9.XI125.NET39_XI9.XI125.MM7_g N_VSS_XI9.XI125.MM7_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.2375e-13 AS=3.225e-13
+ PD=8.95e-07 PS=1.79e-06
mXI9.XI122.MM7 N_XI9.XI122.NET10_XI9.XI122.MM7_d
+ N_XI9.XI122.NET39_XI9.XI122.MM7_g N_VSS_XI9.XI122.MM7_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.2375e-13 AS=3.225e-13
+ PD=8.95e-07 PS=1.79e-06
mXI9.XI114.MM7 N_XI9.XI114.NET10_XI9.XI114.MM7_d
+ N_XI9.XI114.NET39_XI9.XI114.MM7_g N_VSS_XI9.XI114.MM7_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.2375e-13 AS=3.225e-13
+ PD=8.95e-07 PS=1.79e-06
mXI9.XI109.MM7 N_XI9.XI109.NET10_XI9.XI109.MM7_d
+ N_XI9.XI109.NET39_XI9.XI109.MM7_g N_VSS_XI9.XI109.MM7_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.2375e-13 AS=3.225e-13
+ PD=8.95e-07 PS=1.79e-06
mXI9.XI106.MM7 N_XI9.XI106.NET10_XI9.XI106.MM7_d
+ N_XI9.XI106.NET39_XI9.XI106.MM7_g N_VSS_XI9.XI106.MM7_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.2375e-13 AS=3.225e-13
+ PD=8.95e-07 PS=1.79e-06
mXI9.XI101.MM7 N_XI9.XI101.NET10_XI9.XI101.MM7_d
+ N_XI9.XI101.NET39_XI9.XI101.MM7_g N_VSS_XI9.XI101.MM7_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.2375e-13 AS=3.225e-13
+ PD=8.95e-07 PS=1.79e-06
mXI9.XI86.MM7 N_XI9.XI86.NET10_XI9.XI86.MM7_d N_XI9.XI86.NET39_XI9.XI86.MM7_g
+ N_VSS_XI9.XI86.MM7_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.2375e-13 AS=3.225e-13 PD=8.95e-07 PS=1.79e-06
mXI9.XI80.MM7 N_XI9.XI80.NET10_XI9.XI80.MM7_d N_XI9.XI80.NET39_XI9.XI80.MM7_g
+ N_VSS_XI9.XI80.MM7_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.2375e-13 AS=3.225e-13 PD=8.95e-07 PS=1.79e-06
mXI9.XI26.MM7 N_XI9.XI26.NET10_XI9.XI26.MM7_d N_XI9.XI26.NET39_XI9.XI26.MM7_g
+ N_VSS_XI9.XI26.MM7_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.2375e-13 AS=3.225e-13 PD=8.95e-07 PS=1.79e-06
mXI9.XI134.MM6 N_XI9.XI134.NET6_XI9.XI134.MM6_d N_NET241_XI9.XI134.MM6_g
+ N_VSS_XI9.XI134.MM6_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=1.8125e-13 AS=2.575e-13 PD=7.25e-07 PS=1.53e-06
mXI9.XI137.MM2 N_XI9.P15_XI9.XI137.MM2_d N_XI9.XI137.NET43_XI9.XI137.MM2_g
+ N_XI9.XI137.NET10_XI9.XI137.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=4.75e-13 AS=2.2375e-13 PD=1.9e-06 PS=8.95e-07
mXI9.XI140.MM2 N_XI9.P14_XI9.XI140.MM2_d N_XI9.XI140.NET43_XI9.XI140.MM2_g
+ N_XI9.XI140.NET10_XI9.XI140.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=4.75e-13 AS=2.2375e-13 PD=1.9e-06 PS=8.95e-07
mXI9.XI149.MM2 N_XI9.P13_XI9.XI149.MM2_d N_XI9.XI149.NET43_XI9.XI149.MM2_g
+ N_XI9.XI149.NET10_XI9.XI149.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=4.75e-13 AS=2.2375e-13 PD=1.9e-06 PS=8.95e-07
mXI9.XI146.MM2 N_XI9.P12_XI9.XI146.MM2_d N_XI9.XI146.NET43_XI9.XI146.MM2_g
+ N_XI9.XI146.NET10_XI9.XI146.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=4.75e-13 AS=2.2375e-13 PD=1.9e-06 PS=8.95e-07
mXI9.XI143.MM2 N_XI9.P11_XI9.XI143.MM2_d N_XI9.XI143.NET43_XI9.XI143.MM2_g
+ N_XI9.XI143.NET10_XI9.XI143.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=4.75e-13 AS=2.2375e-13 PD=1.9e-06 PS=8.95e-07
mXI9.XI128.MM2 N_XI9.P10_XI9.XI128.MM2_d N_XI9.XI128.NET43_XI9.XI128.MM2_g
+ N_XI9.XI128.NET10_XI9.XI128.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=4.75e-13 AS=2.2375e-13 PD=1.9e-06 PS=8.95e-07
mXI9.XI125.MM2 N_XI9.P9_XI9.XI125.MM2_d N_XI9.XI125.NET43_XI9.XI125.MM2_g
+ N_XI9.XI125.NET10_XI9.XI125.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=4.75e-13 AS=2.2375e-13 PD=1.9e-06 PS=8.95e-07
mXI9.XI122.MM2 N_XI9.P8_XI9.XI122.MM2_d N_XI9.XI122.NET43_XI9.XI122.MM2_g
+ N_XI9.XI122.NET10_XI9.XI122.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=4.75e-13 AS=2.2375e-13 PD=1.9e-06 PS=8.95e-07
mXI9.XI114.MM2 N_XI9.P7_XI9.XI114.MM2_d N_XI9.XI114.NET43_XI9.XI114.MM2_g
+ N_XI9.XI114.NET10_XI9.XI114.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=4.75e-13 AS=2.2375e-13 PD=1.9e-06 PS=8.95e-07
mXI9.XI109.MM2 N_XI9.P6_XI9.XI109.MM2_d N_XI9.XI109.NET43_XI9.XI109.MM2_g
+ N_XI9.XI109.NET10_XI9.XI109.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=4.75e-13 AS=2.2375e-13 PD=1.9e-06 PS=8.95e-07
mXI9.XI106.MM2 N_XI9.P5_XI9.XI106.MM2_d N_XI9.XI106.NET43_XI9.XI106.MM2_g
+ N_XI9.XI106.NET10_XI9.XI106.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=4.75e-13 AS=2.2375e-13 PD=1.9e-06 PS=8.95e-07
mXI9.XI101.MM2 N_XI9.P4_XI9.XI101.MM2_d N_XI9.XI101.NET43_XI9.XI101.MM2_g
+ N_XI9.XI101.NET10_XI9.XI101.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=4.75e-13 AS=2.2375e-13 PD=1.9e-06 PS=8.95e-07
mXI9.XI86.MM2 N_XI9.P3_XI9.XI86.MM2_d N_XI9.XI86.NET43_XI9.XI86.MM2_g
+ N_XI9.XI86.NET10_XI9.XI86.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=4.75e-13 AS=2.2375e-13 PD=1.9e-06 PS=8.95e-07
mXI9.XI80.MM2 N_XI9.P2_XI9.XI80.MM2_d N_XI9.XI80.NET43_XI9.XI80.MM2_g
+ N_XI9.XI80.NET10_XI9.XI80.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=4.75e-13 AS=2.2375e-13 PD=1.9e-06 PS=8.95e-07
mXI9.XI26.MM2 N_XI9.P1_XI9.XI26.MM2_d N_XI9.XI26.NET43_XI9.XI26.MM2_g
+ N_XI9.XI26.NET10_XI9.XI26.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=4.75e-13 AS=2.2375e-13 PD=1.9e-06 PS=8.95e-07
mXI9.XI134.XI9.MM2 N_XI9.XI134.NET43_XI9.XI134.XI9.MM2_d
+ N_ACC15_XI9.XI134.XI9.MM2_g N_VSS_XI9.XI134.XI9.MM2_s N_VSS_XI10.XI0.XI0.MM2_b
+ N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9.XI137.MM0 N_XI9.P15_XI9.XI137.MM0_d N_ACC14_XI9.XI137.MM0_g
+ N_XI9.XI137.NET6_XI9.XI137.MM0_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=4.75e-13 AS=1.8125e-13 PD=1.9e-06 PS=7.25e-07
mXI9.XI140.MM0 N_XI9.P14_XI9.XI140.MM0_d N_ACC13_XI9.XI140.MM0_g
+ N_XI9.XI140.NET6_XI9.XI140.MM0_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=4.75e-13 AS=1.8125e-13 PD=1.9e-06 PS=7.25e-07
mXI9.XI149.MM0 N_XI9.P13_XI9.XI149.MM0_d N_ACC12_XI9.XI149.MM0_g
+ N_XI9.XI149.NET6_XI9.XI149.MM0_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=4.75e-13 AS=1.8125e-13 PD=1.9e-06 PS=7.25e-07
mXI9.XI146.MM0 N_XI9.P12_XI9.XI146.MM0_d N_ACC11_XI9.XI146.MM0_g
+ N_XI9.XI146.NET6_XI9.XI146.MM0_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=4.75e-13 AS=1.8125e-13 PD=1.9e-06 PS=7.25e-07
mXI9.XI143.MM0 N_XI9.P11_XI9.XI143.MM0_d N_ACC10_XI9.XI143.MM0_g
+ N_XI9.XI143.NET6_XI9.XI143.MM0_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=4.75e-13 AS=1.8125e-13 PD=1.9e-06 PS=7.25e-07
mXI9.XI128.MM0 N_XI9.P10_XI9.XI128.MM0_d N_ACC9_XI9.XI128.MM0_g
+ N_XI9.XI128.NET6_XI9.XI128.MM0_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=4.75e-13 AS=1.8125e-13 PD=1.9e-06 PS=7.25e-07
mXI9.XI125.MM0 N_XI9.P9_XI9.XI125.MM0_d N_ACC8_XI9.XI125.MM0_g
+ N_XI9.XI125.NET6_XI9.XI125.MM0_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=4.75e-13 AS=1.8125e-13 PD=1.9e-06 PS=7.25e-07
mXI9.XI122.MM0 N_XI9.P8_XI9.XI122.MM0_d N_ACC7_XI9.XI122.MM0_g
+ N_XI9.XI122.NET6_XI9.XI122.MM0_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=4.75e-13 AS=1.8125e-13 PD=1.9e-06 PS=7.25e-07
mXI9.XI114.MM0 N_XI9.P7_XI9.XI114.MM0_d N_ACC6_XI9.XI114.MM0_g
+ N_XI9.XI114.NET6_XI9.XI114.MM0_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=4.75e-13 AS=1.8125e-13 PD=1.9e-06 PS=7.25e-07
mXI9.XI109.MM0 N_XI9.P6_XI9.XI109.MM0_d N_ACC5_XI9.XI109.MM0_g
+ N_XI9.XI109.NET6_XI9.XI109.MM0_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=4.75e-13 AS=1.8125e-13 PD=1.9e-06 PS=7.25e-07
mXI9.XI106.MM0 N_XI9.P5_XI9.XI106.MM0_d N_ACC4_XI9.XI106.MM0_g
+ N_XI9.XI106.NET6_XI9.XI106.MM0_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=4.75e-13 AS=1.8125e-13 PD=1.9e-06 PS=7.25e-07
mXI9.XI101.MM0 N_XI9.P4_XI9.XI101.MM0_d N_ACC3_XI9.XI101.MM0_g
+ N_XI9.XI101.NET6_XI9.XI101.MM0_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=4.75e-13 AS=1.8125e-13 PD=1.9e-06 PS=7.25e-07
mXI9.XI86.MM0 N_XI9.P3_XI9.XI86.MM0_d N_ACC2_XI9.XI86.MM0_g
+ N_XI9.XI86.NET6_XI9.XI86.MM0_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=4.75e-13 AS=1.8125e-13 PD=1.9e-06 PS=7.25e-07
mXI9.XI80.MM0 N_XI9.P2_XI9.XI80.MM0_d N_ACC1_XI9.XI80.MM0_g
+ N_XI9.XI80.NET6_XI9.XI80.MM0_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=4.75e-13 AS=1.8125e-13 PD=1.9e-06 PS=7.25e-07
mXI9.XI26.MM0 N_XI9.P1_XI9.XI26.MM0_d N_ACC0_XI9.XI26.MM0_g
+ N_XI9.XI26.NET6_XI9.XI26.MM0_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=4.75e-13 AS=1.8125e-13 PD=1.9e-06 PS=7.25e-07
mXI9.XI137.MM6 N_XI9.XI137.NET6_XI9.XI137.MM6_d N_NET242_XI9.XI137.MM6_g
+ N_VSS_XI9.XI137.MM6_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=1.8125e-13 AS=2.575e-13 PD=7.25e-07 PS=1.53e-06
mXI9.XI140.MM6 N_XI9.XI140.NET6_XI9.XI140.MM6_d N_NET243_XI9.XI140.MM6_g
+ N_VSS_XI9.XI140.MM6_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=1.8125e-13 AS=2.575e-13 PD=7.25e-07 PS=1.53e-06
mXI9.XI149.MM6 N_XI9.XI149.NET6_XI9.XI149.MM6_d N_NET244_XI9.XI149.MM6_g
+ N_VSS_XI9.XI149.MM6_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=1.8125e-13 AS=2.575e-13 PD=7.25e-07 PS=1.53e-06
mXI9.XI146.MM6 N_XI9.XI146.NET6_XI9.XI146.MM6_d N_NET245_XI9.XI146.MM6_g
+ N_VSS_XI9.XI146.MM6_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=1.8125e-13 AS=2.575e-13 PD=7.25e-07 PS=1.53e-06
mXI9.XI143.MM6 N_XI9.XI143.NET6_XI9.XI143.MM6_d N_NET246_XI9.XI143.MM6_g
+ N_VSS_XI9.XI143.MM6_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=1.8125e-13 AS=2.575e-13 PD=7.25e-07 PS=1.53e-06
mXI9.XI128.MM6 N_XI9.XI128.NET6_XI9.XI128.MM6_d N_NET247_XI9.XI128.MM6_g
+ N_VSS_XI9.XI128.MM6_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=1.8125e-13 AS=2.575e-13 PD=7.25e-07 PS=1.53e-06
mXI9.XI125.MM6 N_XI9.XI125.NET6_XI9.XI125.MM6_d N_NET248_XI9.XI125.MM6_g
+ N_VSS_XI9.XI125.MM6_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=1.8125e-13 AS=2.575e-13 PD=7.25e-07 PS=1.53e-06
mXI9.XI122.MM6 N_XI9.XI122.NET6_XI9.XI122.MM6_d N_NET249_XI9.XI122.MM6_g
+ N_VSS_XI9.XI122.MM6_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=1.8125e-13 AS=2.575e-13 PD=7.25e-07 PS=1.53e-06
mXI9.XI114.MM6 N_XI9.XI114.NET6_XI9.XI114.MM6_d N_NET250_XI9.XI114.MM6_g
+ N_VSS_XI9.XI114.MM6_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=1.8125e-13 AS=2.575e-13 PD=7.25e-07 PS=1.53e-06
mXI9.XI109.MM6 N_XI9.XI109.NET6_XI9.XI109.MM6_d N_NET251_XI9.XI109.MM6_g
+ N_VSS_XI9.XI109.MM6_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=1.8125e-13 AS=2.575e-13 PD=7.25e-07 PS=1.53e-06
mXI9.XI106.MM6 N_XI9.XI106.NET6_XI9.XI106.MM6_d N_NET252_XI9.XI106.MM6_g
+ N_VSS_XI9.XI106.MM6_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=1.8125e-13 AS=2.575e-13 PD=7.25e-07 PS=1.53e-06
mXI9.XI101.MM6 N_XI9.XI101.NET6_XI9.XI101.MM6_d N_NET253_XI9.XI101.MM6_g
+ N_VSS_XI9.XI101.MM6_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=1.8125e-13 AS=2.575e-13 PD=7.25e-07 PS=1.53e-06
mXI9.XI86.MM6 N_XI9.XI86.NET6_XI9.XI86.MM6_d N_NET254_XI9.XI86.MM6_g
+ N_VSS_XI9.XI86.MM6_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=1.8125e-13 AS=2.575e-13 PD=7.25e-07 PS=1.53e-06
mXI9.XI80.MM6 N_XI9.XI80.NET6_XI9.XI80.MM6_d N_NET255_XI9.XI80.MM6_g
+ N_VSS_XI9.XI80.MM6_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=1.8125e-13 AS=2.575e-13 PD=7.25e-07 PS=1.53e-06
mXI9.XI26.MM6 N_XI9.XI26.NET6_XI9.XI26.MM6_d N_NET256_XI9.XI26.MM6_g
+ N_VSS_XI9.XI26.MM6_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=1.8125e-13 AS=2.575e-13 PD=7.25e-07 PS=1.53e-06
mXI9.XI137.XI9.MM2 N_XI9.XI137.NET43_XI9.XI137.XI9.MM2_d
+ N_ACC14_XI9.XI137.XI9.MM2_g N_VSS_XI9.XI137.XI9.MM2_s N_VSS_XI10.XI0.XI0.MM2_b
+ N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9.XI140.XI9.MM2 N_XI9.XI140.NET43_XI9.XI140.XI9.MM2_d
+ N_ACC13_XI9.XI140.XI9.MM2_g N_VSS_XI9.XI140.XI9.MM2_s N_VSS_XI10.XI0.XI0.MM2_b
+ N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9.XI149.XI9.MM2 N_XI9.XI149.NET43_XI9.XI149.XI9.MM2_d
+ N_ACC12_XI9.XI149.XI9.MM2_g N_VSS_XI9.XI149.XI9.MM2_s N_VSS_XI10.XI0.XI0.MM2_b
+ N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9.XI146.XI9.MM2 N_XI9.XI146.NET43_XI9.XI146.XI9.MM2_d
+ N_ACC11_XI9.XI146.XI9.MM2_g N_VSS_XI9.XI146.XI9.MM2_s N_VSS_XI10.XI0.XI0.MM2_b
+ N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9.XI143.XI9.MM2 N_XI9.XI143.NET43_XI9.XI143.XI9.MM2_d
+ N_ACC10_XI9.XI143.XI9.MM2_g N_VSS_XI9.XI143.XI9.MM2_s N_VSS_XI10.XI0.XI0.MM2_b
+ N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9.XI128.XI9.MM2 N_XI9.XI128.NET43_XI9.XI128.XI9.MM2_d
+ N_ACC9_XI9.XI128.XI9.MM2_g N_VSS_XI9.XI128.XI9.MM2_s N_VSS_XI10.XI0.XI0.MM2_b
+ N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9.XI125.XI9.MM2 N_XI9.XI125.NET43_XI9.XI125.XI9.MM2_d
+ N_ACC8_XI9.XI125.XI9.MM2_g N_VSS_XI9.XI125.XI9.MM2_s N_VSS_XI10.XI0.XI0.MM2_b
+ N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9.XI122.XI9.MM2 N_XI9.XI122.NET43_XI9.XI122.XI9.MM2_d
+ N_ACC7_XI9.XI122.XI9.MM2_g N_VSS_XI9.XI122.XI9.MM2_s N_VSS_XI10.XI0.XI0.MM2_b
+ N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9.XI114.XI9.MM2 N_XI9.XI114.NET43_XI9.XI114.XI9.MM2_d
+ N_ACC6_XI9.XI114.XI9.MM2_g N_VSS_XI9.XI114.XI9.MM2_s N_VSS_XI10.XI0.XI0.MM2_b
+ N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9.XI109.XI9.MM2 N_XI9.XI109.NET43_XI9.XI109.XI9.MM2_d
+ N_ACC5_XI9.XI109.XI9.MM2_g N_VSS_XI9.XI109.XI9.MM2_s N_VSS_XI10.XI0.XI0.MM2_b
+ N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9.XI106.XI9.MM2 N_XI9.XI106.NET43_XI9.XI106.XI9.MM2_d
+ N_ACC4_XI9.XI106.XI9.MM2_g N_VSS_XI9.XI106.XI9.MM2_s N_VSS_XI10.XI0.XI0.MM2_b
+ N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9.XI101.XI9.MM2 N_XI9.XI101.NET43_XI9.XI101.XI9.MM2_d
+ N_ACC3_XI9.XI101.XI9.MM2_g N_VSS_XI9.XI101.XI9.MM2_s N_VSS_XI10.XI0.XI0.MM2_b
+ N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9.XI86.XI9.MM2 N_XI9.XI86.NET43_XI9.XI86.XI9.MM2_d N_ACC2_XI9.XI86.XI9.MM2_g
+ N_VSS_XI9.XI86.XI9.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9.XI80.XI9.MM2 N_XI9.XI80.NET43_XI9.XI80.XI9.MM2_d N_ACC1_XI9.XI80.XI9.MM2_g
+ N_VSS_XI9.XI80.XI9.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9.XI26.XI9.MM2 N_XI9.XI26.NET43_XI9.XI26.XI9.MM2_d N_ACC0_XI9.XI26.XI9.MM2_g
+ N_VSS_XI9.XI26.XI9.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9.XI168.XI1.XI1.MM0 N_XI9.XI168.XI1.XI1.NET036_XI9.XI168.XI1.XI1.MM0_d
+ N_XI9.NET138_XI9.XI168.XI1.XI1.MM0_g N_VSS_XI9.XI168.XI1.XI1.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.85e-13 AS=2.45e-13
+ PD=7.4e-07 PS=1.48e-06
mXI9.XI167.XI1.XI1.MM0 N_XI9.XI167.XI1.XI1.NET036_XI9.XI167.XI1.XI1.MM0_d
+ N_XI9.NET208_XI9.XI167.XI1.XI1.MM0_g N_VSS_XI9.XI167.XI1.XI1.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.85e-13 AS=2.45e-13
+ PD=7.4e-07 PS=1.48e-06
mXI9.XI166.XI1.XI1.MM0 N_XI9.XI166.XI1.XI1.NET036_XI9.XI166.XI1.XI1.MM0_d
+ N_XI9.NET202_XI9.XI166.XI1.XI1.MM0_g N_VSS_XI9.XI166.XI1.XI1.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.85e-13 AS=2.45e-13
+ PD=7.4e-07 PS=1.48e-06
mXI9.XI165.XI1.XI1.MM0 N_XI9.XI165.XI1.XI1.NET036_XI9.XI165.XI1.XI1.MM0_d
+ N_XI9.NET198_XI9.XI165.XI1.XI1.MM0_g N_VSS_XI9.XI165.XI1.XI1.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.85e-13 AS=2.45e-13
+ PD=7.4e-07 PS=1.48e-06
mXI9.XI159.XI1.XI1.MM0 N_XI9.XI159.XI1.XI1.NET036_XI9.XI159.XI1.XI1.MM0_d
+ N_XI9.NET102_XI9.XI159.XI1.XI1.MM0_g N_VSS_XI9.XI159.XI1.XI1.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.85e-13 AS=2.45e-13
+ PD=7.4e-07 PS=1.48e-06
mXI9.XI160.XI1.XI1.MM0 N_XI9.XI160.XI1.XI1.NET036_XI9.XI160.XI1.XI1.MM0_d
+ N_XI9.NET108_XI9.XI160.XI1.XI1.MM0_g N_VSS_XI9.XI160.XI1.XI1.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.85e-13 AS=2.45e-13
+ PD=7.4e-07 PS=1.48e-06
mXI9.XI161.XI1.XI1.MM0 N_XI9.XI161.XI1.XI1.NET036_XI9.XI161.XI1.XI1.MM0_d
+ N_XI9.NET96_XI9.XI161.XI1.XI1.MM0_g N_VSS_XI9.XI161.XI1.XI1.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.85e-13 AS=2.45e-13
+ PD=7.4e-07 PS=1.48e-06
mXI9.XI162.XI1.XI1.MM0 N_XI9.XI162.XI1.XI1.NET036_XI9.XI162.XI1.XI1.MM0_d
+ N_XI9.NET153_XI9.XI162.XI1.XI1.MM0_g N_VSS_XI9.XI162.XI1.XI1.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.85e-13 AS=2.45e-13
+ PD=7.4e-07 PS=1.48e-06
mXI9.XI121.XI1.XI1.MM0 N_XI9.XI121.XI1.XI1.NET036_XI9.XI121.XI1.XI1.MM0_d
+ N_XI9.NET54_XI9.XI121.XI1.XI1.MM0_g N_VSS_XI9.XI121.XI1.XI1.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.85e-13 AS=2.45e-13
+ PD=7.4e-07 PS=1.48e-06
mXI9.XI120.XI1.XI1.MM0 N_XI9.XI120.XI1.XI1.NET036_XI9.XI120.XI1.XI1.MM0_d
+ N_XI9.NET66_XI9.XI120.XI1.XI1.MM0_g N_VSS_XI9.XI120.XI1.XI1.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.85e-13 AS=2.45e-13
+ PD=7.4e-07 PS=1.48e-06
mXI9.XI119.XI1.XI1.MM0 N_XI9.XI119.XI1.XI1.NET036_XI9.XI119.XI1.XI1.MM0_d
+ N_XI9.NET72_XI9.XI119.XI1.XI1.MM0_g N_VSS_XI9.XI119.XI1.XI1.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.85e-13 AS=2.45e-13
+ PD=7.4e-07 PS=1.48e-06
mXI9.XI118.XI1.XI1.MM0 N_XI9.XI118.XI1.XI1.NET036_XI9.XI118.XI1.XI1.MM0_d
+ N_XI9.NET60_XI9.XI118.XI1.XI1.MM0_g N_VSS_XI9.XI118.XI1.XI1.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.85e-13 AS=2.45e-13
+ PD=7.4e-07 PS=1.48e-06
mXI9.XI91.XI1.XI1.MM0 N_XI9.XI91.XI1.XI1.NET036_XI9.XI91.XI1.XI1.MM0_d
+ N_XI9.NET183_XI9.XI91.XI1.XI1.MM0_g N_VSS_XI9.XI91.XI1.XI1.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.85e-13 AS=2.45e-13
+ PD=7.4e-07 PS=1.48e-06
mXI9.XI90.XI1.XI1.MM0 N_XI9.XI90.XI1.XI1.NET036_XI9.XI90.XI1.XI1.MM0_d
+ N_XI9.NET178_XI9.XI90.XI1.XI1.MM0_g N_VSS_XI9.XI90.XI1.XI1.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.85e-13 AS=2.45e-13
+ PD=7.4e-07 PS=1.48e-06
mXI9.XI89.XI1.XI1.MM0 N_XI9.XI89.XI1.XI1.NET036_XI9.XI89.XI1.XI1.MM0_d
+ N_CIN1_XI9.XI89.XI1.XI1.MM0_g N_VSS_XI9.XI89.XI1.XI1.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.85e-13 AS=2.45e-13
+ PD=7.4e-07 PS=1.48e-06
mXI9.XI168.XI1.XI1.MM2 N_XI9.XI168.XI1.NET6_XI9.XI168.XI1.XI1.MM2_d
+ N_XI9.P15_XI9.XI168.XI1.XI1.MM2_g
+ N_XI9.XI168.XI1.XI1.NET036_XI9.XI168.XI1.XI1.MM2_s N_VSS_XI10.XI0.XI0.MM2_b
+ N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=1.85e-13 PD=1.52e-06 PS=7.4e-07
mXI9.XI167.XI1.XI1.MM2 N_XI9.XI167.XI1.NET6_XI9.XI167.XI1.XI1.MM2_d
+ N_XI9.P14_XI9.XI167.XI1.XI1.MM2_g
+ N_XI9.XI167.XI1.XI1.NET036_XI9.XI167.XI1.XI1.MM2_s N_VSS_XI10.XI0.XI0.MM2_b
+ N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=1.85e-13 PD=1.52e-06 PS=7.4e-07
mXI9.XI166.XI1.XI1.MM2 N_XI9.XI166.XI1.NET6_XI9.XI166.XI1.XI1.MM2_d
+ N_XI9.P13_XI9.XI166.XI1.XI1.MM2_g
+ N_XI9.XI166.XI1.XI1.NET036_XI9.XI166.XI1.XI1.MM2_s N_VSS_XI10.XI0.XI0.MM2_b
+ N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=1.85e-13 PD=1.52e-06 PS=7.4e-07
mXI9.XI165.XI1.XI1.MM2 N_XI9.XI165.XI1.NET6_XI9.XI165.XI1.XI1.MM2_d
+ N_XI9.P12_XI9.XI165.XI1.XI1.MM2_g
+ N_XI9.XI165.XI1.XI1.NET036_XI9.XI165.XI1.XI1.MM2_s N_VSS_XI10.XI0.XI0.MM2_b
+ N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=1.85e-13 PD=1.52e-06 PS=7.4e-07
mXI9.XI159.XI1.XI1.MM2 N_XI9.XI159.XI1.NET6_XI9.XI159.XI1.XI1.MM2_d
+ N_XI9.P11_XI9.XI159.XI1.XI1.MM2_g
+ N_XI9.XI159.XI1.XI1.NET036_XI9.XI159.XI1.XI1.MM2_s N_VSS_XI10.XI0.XI0.MM2_b
+ N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=1.85e-13 PD=1.52e-06 PS=7.4e-07
mXI9.XI160.XI1.XI1.MM2 N_XI9.XI160.XI1.NET6_XI9.XI160.XI1.XI1.MM2_d
+ N_XI9.P10_XI9.XI160.XI1.XI1.MM2_g
+ N_XI9.XI160.XI1.XI1.NET036_XI9.XI160.XI1.XI1.MM2_s N_VSS_XI10.XI0.XI0.MM2_b
+ N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=1.85e-13 PD=1.52e-06 PS=7.4e-07
mXI9.XI161.XI1.XI1.MM2 N_XI9.XI161.XI1.NET6_XI9.XI161.XI1.XI1.MM2_d
+ N_XI9.P9_XI9.XI161.XI1.XI1.MM2_g
+ N_XI9.XI161.XI1.XI1.NET036_XI9.XI161.XI1.XI1.MM2_s N_VSS_XI10.XI0.XI0.MM2_b
+ N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=1.85e-13 PD=1.52e-06 PS=7.4e-07
mXI9.XI162.XI1.XI1.MM2 N_XI9.XI162.XI1.NET6_XI9.XI162.XI1.XI1.MM2_d
+ N_XI9.P8_XI9.XI162.XI1.XI1.MM2_g
+ N_XI9.XI162.XI1.XI1.NET036_XI9.XI162.XI1.XI1.MM2_s N_VSS_XI10.XI0.XI0.MM2_b
+ N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=1.85e-13 PD=1.52e-06 PS=7.4e-07
mXI9.XI121.XI1.XI1.MM2 N_XI9.XI121.XI1.NET6_XI9.XI121.XI1.XI1.MM2_d
+ N_XI9.P7_XI9.XI121.XI1.XI1.MM2_g
+ N_XI9.XI121.XI1.XI1.NET036_XI9.XI121.XI1.XI1.MM2_s N_VSS_XI10.XI0.XI0.MM2_b
+ N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=1.85e-13 PD=1.52e-06 PS=7.4e-07
mXI9.XI120.XI1.XI1.MM2 N_XI9.XI120.XI1.NET6_XI9.XI120.XI1.XI1.MM2_d
+ N_XI9.P6_XI9.XI120.XI1.XI1.MM2_g
+ N_XI9.XI120.XI1.XI1.NET036_XI9.XI120.XI1.XI1.MM2_s N_VSS_XI10.XI0.XI0.MM2_b
+ N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=1.85e-13 PD=1.52e-06 PS=7.4e-07
mXI9.XI119.XI1.XI1.MM2 N_XI9.XI119.XI1.NET6_XI9.XI119.XI1.XI1.MM2_d
+ N_XI9.P5_XI9.XI119.XI1.XI1.MM2_g
+ N_XI9.XI119.XI1.XI1.NET036_XI9.XI119.XI1.XI1.MM2_s N_VSS_XI10.XI0.XI0.MM2_b
+ N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=1.85e-13 PD=1.52e-06 PS=7.4e-07
mXI9.XI118.XI1.XI1.MM2 N_XI9.XI118.XI1.NET6_XI9.XI118.XI1.XI1.MM2_d
+ N_XI9.P4_XI9.XI118.XI1.XI1.MM2_g
+ N_XI9.XI118.XI1.XI1.NET036_XI9.XI118.XI1.XI1.MM2_s N_VSS_XI10.XI0.XI0.MM2_b
+ N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=1.85e-13 PD=1.52e-06 PS=7.4e-07
mXI9.XI91.XI1.XI1.MM2 N_XI9.XI91.XI1.NET6_XI9.XI91.XI1.XI1.MM2_d
+ N_XI9.P3_XI9.XI91.XI1.XI1.MM2_g
+ N_XI9.XI91.XI1.XI1.NET036_XI9.XI91.XI1.XI1.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18
+ L=1.8e-07 W=5e-07 AD=2.55e-13 AS=1.85e-13 PD=1.52e-06 PS=7.4e-07
mXI9.XI90.XI1.XI1.MM2 N_XI9.XI90.XI1.NET6_XI9.XI90.XI1.XI1.MM2_d
+ N_XI9.P2_XI9.XI90.XI1.XI1.MM2_g
+ N_XI9.XI90.XI1.XI1.NET036_XI9.XI90.XI1.XI1.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18
+ L=1.8e-07 W=5e-07 AD=2.55e-13 AS=1.85e-13 PD=1.52e-06 PS=7.4e-07
mXI9.XI89.XI1.XI1.MM2 N_XI9.XI89.XI1.NET6_XI9.XI89.XI1.XI1.MM2_d
+ N_XI9.P1_XI9.XI89.XI1.XI1.MM2_g
+ N_XI9.XI89.XI1.XI1.NET036_XI9.XI89.XI1.XI1.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18
+ L=1.8e-07 W=5e-07 AD=2.55e-13 AS=1.85e-13 PD=1.52e-06 PS=7.4e-07
mXI9.XI168.XI1.XI0.MM2 N_XI9.XI168.NET13_XI9.XI168.XI1.XI0.MM2_d
+ N_XI9.XI168.XI1.NET6_XI9.XI168.XI1.XI0.MM2_g N_VSS_XI9.XI168.XI1.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI9.XI167.XI1.XI0.MM2 N_XI9.XI167.NET13_XI9.XI167.XI1.XI0.MM2_d
+ N_XI9.XI167.XI1.NET6_XI9.XI167.XI1.XI0.MM2_g N_VSS_XI9.XI167.XI1.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI9.XI166.XI1.XI0.MM2 N_XI9.XI166.NET13_XI9.XI166.XI1.XI0.MM2_d
+ N_XI9.XI166.XI1.NET6_XI9.XI166.XI1.XI0.MM2_g N_VSS_XI9.XI166.XI1.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI9.XI165.XI1.XI0.MM2 N_XI9.XI165.NET13_XI9.XI165.XI1.XI0.MM2_d
+ N_XI9.XI165.XI1.NET6_XI9.XI165.XI1.XI0.MM2_g N_VSS_XI9.XI165.XI1.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI9.XI159.XI1.XI0.MM2 N_XI9.XI159.NET13_XI9.XI159.XI1.XI0.MM2_d
+ N_XI9.XI159.XI1.NET6_XI9.XI159.XI1.XI0.MM2_g N_VSS_XI9.XI159.XI1.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI9.XI160.XI1.XI0.MM2 N_XI9.XI160.NET13_XI9.XI160.XI1.XI0.MM2_d
+ N_XI9.XI160.XI1.NET6_XI9.XI160.XI1.XI0.MM2_g N_VSS_XI9.XI160.XI1.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI9.XI161.XI1.XI0.MM2 N_XI9.XI161.NET13_XI9.XI161.XI1.XI0.MM2_d
+ N_XI9.XI161.XI1.NET6_XI9.XI161.XI1.XI0.MM2_g N_VSS_XI9.XI161.XI1.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI9.XI162.XI1.XI0.MM2 N_XI9.XI162.NET13_XI9.XI162.XI1.XI0.MM2_d
+ N_XI9.XI162.XI1.NET6_XI9.XI162.XI1.XI0.MM2_g N_VSS_XI9.XI162.XI1.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI9.XI121.XI1.XI0.MM2 N_XI9.XI121.NET13_XI9.XI121.XI1.XI0.MM2_d
+ N_XI9.XI121.XI1.NET6_XI9.XI121.XI1.XI0.MM2_g N_VSS_XI9.XI121.XI1.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI9.XI120.XI1.XI0.MM2 N_XI9.XI120.NET13_XI9.XI120.XI1.XI0.MM2_d
+ N_XI9.XI120.XI1.NET6_XI9.XI120.XI1.XI0.MM2_g N_VSS_XI9.XI120.XI1.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI9.XI119.XI1.XI0.MM2 N_XI9.XI119.NET13_XI9.XI119.XI1.XI0.MM2_d
+ N_XI9.XI119.XI1.NET6_XI9.XI119.XI1.XI0.MM2_g N_VSS_XI9.XI119.XI1.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI9.XI118.XI1.XI0.MM2 N_XI9.XI118.NET13_XI9.XI118.XI1.XI0.MM2_d
+ N_XI9.XI118.XI1.NET6_XI9.XI118.XI1.XI0.MM2_g N_VSS_XI9.XI118.XI1.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI9.XI91.XI1.XI0.MM2 N_XI9.XI91.NET13_XI9.XI91.XI1.XI0.MM2_d
+ N_XI9.XI91.XI1.NET6_XI9.XI91.XI1.XI0.MM2_g N_VSS_XI9.XI91.XI1.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI9.XI90.XI1.XI0.MM2 N_XI9.XI90.NET13_XI9.XI90.XI1.XI0.MM2_d
+ N_XI9.XI90.XI1.NET6_XI9.XI90.XI1.XI0.MM2_g N_VSS_XI9.XI90.XI1.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI9.XI89.XI1.XI0.MM2 N_XI9.XI89.NET13_XI9.XI89.XI1.XI0.MM2_d
+ N_XI9.XI89.XI1.NET6_XI9.XI89.XI1.XI0.MM2_g N_VSS_XI9.XI89.XI1.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI9.XI168.XI0.XI0.MM0 N_XI9.XI168.XI0.NET12_XI9.XI168.XI0.XI0.MM0_d
+ N_XI9.XI168.NET13_XI9.XI168.XI0.XI0.MM0_g N_VSS_XI9.XI168.XI0.XI0.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.375e-13 AS=2.45e-13
+ PD=5.5e-07 PS=1.48e-06
mXI9.XI167.XI0.XI0.MM0 N_XI9.XI167.XI0.NET12_XI9.XI167.XI0.XI0.MM0_d
+ N_XI9.XI167.NET13_XI9.XI167.XI0.XI0.MM0_g N_VSS_XI9.XI167.XI0.XI0.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.375e-13 AS=2.45e-13
+ PD=5.5e-07 PS=1.48e-06
mXI9.XI166.XI0.XI0.MM0 N_XI9.XI166.XI0.NET12_XI9.XI166.XI0.XI0.MM0_d
+ N_XI9.XI166.NET13_XI9.XI166.XI0.XI0.MM0_g N_VSS_XI9.XI166.XI0.XI0.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.375e-13 AS=2.45e-13
+ PD=5.5e-07 PS=1.48e-06
mXI9.XI165.XI0.XI0.MM0 N_XI9.XI165.XI0.NET12_XI9.XI165.XI0.XI0.MM0_d
+ N_XI9.XI165.NET13_XI9.XI165.XI0.XI0.MM0_g N_VSS_XI9.XI165.XI0.XI0.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.375e-13 AS=2.45e-13
+ PD=5.5e-07 PS=1.48e-06
mXI9.XI159.XI0.XI0.MM0 N_XI9.XI159.XI0.NET12_XI9.XI159.XI0.XI0.MM0_d
+ N_XI9.XI159.NET13_XI9.XI159.XI0.XI0.MM0_g N_VSS_XI9.XI159.XI0.XI0.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.375e-13 AS=2.45e-13
+ PD=5.5e-07 PS=1.48e-06
mXI9.XI160.XI0.XI0.MM0 N_XI9.XI160.XI0.NET12_XI9.XI160.XI0.XI0.MM0_d
+ N_XI9.XI160.NET13_XI9.XI160.XI0.XI0.MM0_g N_VSS_XI9.XI160.XI0.XI0.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.375e-13 AS=2.45e-13
+ PD=5.5e-07 PS=1.48e-06
mXI9.XI161.XI0.XI0.MM0 N_XI9.XI161.XI0.NET12_XI9.XI161.XI0.XI0.MM0_d
+ N_XI9.XI161.NET13_XI9.XI161.XI0.XI0.MM0_g N_VSS_XI9.XI161.XI0.XI0.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.375e-13 AS=2.45e-13
+ PD=5.5e-07 PS=1.48e-06
mXI9.XI162.XI0.XI0.MM0 N_XI9.XI162.XI0.NET12_XI9.XI162.XI0.XI0.MM0_d
+ N_XI9.XI162.NET13_XI9.XI162.XI0.XI0.MM0_g N_VSS_XI9.XI162.XI0.XI0.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.375e-13 AS=2.45e-13
+ PD=5.5e-07 PS=1.48e-06
mXI9.XI121.XI0.XI0.MM0 N_XI9.XI121.XI0.NET12_XI9.XI121.XI0.XI0.MM0_d
+ N_XI9.XI121.NET13_XI9.XI121.XI0.XI0.MM0_g N_VSS_XI9.XI121.XI0.XI0.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.375e-13 AS=2.45e-13
+ PD=5.5e-07 PS=1.48e-06
mXI9.XI120.XI0.XI0.MM0 N_XI9.XI120.XI0.NET12_XI9.XI120.XI0.XI0.MM0_d
+ N_XI9.XI120.NET13_XI9.XI120.XI0.XI0.MM0_g N_VSS_XI9.XI120.XI0.XI0.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.375e-13 AS=2.45e-13
+ PD=5.5e-07 PS=1.48e-06
mXI9.XI119.XI0.XI0.MM0 N_XI9.XI119.XI0.NET12_XI9.XI119.XI0.XI0.MM0_d
+ N_XI9.XI119.NET13_XI9.XI119.XI0.XI0.MM0_g N_VSS_XI9.XI119.XI0.XI0.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.375e-13 AS=2.45e-13
+ PD=5.5e-07 PS=1.48e-06
mXI9.XI118.XI0.XI0.MM0 N_XI9.XI118.XI0.NET12_XI9.XI118.XI0.XI0.MM0_d
+ N_XI9.XI118.NET13_XI9.XI118.XI0.XI0.MM0_g N_VSS_XI9.XI118.XI0.XI0.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.375e-13 AS=2.45e-13
+ PD=5.5e-07 PS=1.48e-06
mXI9.XI91.XI0.XI0.MM0 N_XI9.XI91.XI0.NET12_XI9.XI91.XI0.XI0.MM0_d
+ N_XI9.XI91.NET13_XI9.XI91.XI0.XI0.MM0_g N_VSS_XI9.XI91.XI0.XI0.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.375e-13 AS=2.45e-13
+ PD=5.5e-07 PS=1.48e-06
mXI9.XI90.XI0.XI0.MM0 N_XI9.XI90.XI0.NET12_XI9.XI90.XI0.XI0.MM0_d
+ N_XI9.XI90.NET13_XI9.XI90.XI0.XI0.MM0_g N_VSS_XI9.XI90.XI0.XI0.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.375e-13 AS=2.45e-13
+ PD=5.5e-07 PS=1.48e-06
mXI9.XI89.XI0.XI0.MM0 N_XI9.XI89.XI0.NET12_XI9.XI89.XI0.XI0.MM0_d
+ N_XI9.XI89.NET13_XI9.XI89.XI0.XI0.MM0_g N_VSS_XI9.XI89.XI0.XI0.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.375e-13 AS=2.45e-13
+ PD=5.5e-07 PS=1.48e-06
mXI9.XI168.XI0.XI0.MM2 N_XI9.XI168.XI0.NET12_XI9.XI168.XI0.XI0.MM2_d
+ N_XI9.G15_XI9.XI168.XI0.XI0.MM2_g N_VSS_XI9.XI168.XI0.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.375e-13 AS=2.55e-13
+ PD=5.5e-07 PS=1.52e-06
mXI9.XI167.XI0.XI0.MM2 N_XI9.XI167.XI0.NET12_XI9.XI167.XI0.XI0.MM2_d
+ N_XI9.G14_XI9.XI167.XI0.XI0.MM2_g N_VSS_XI9.XI167.XI0.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.375e-13 AS=2.55e-13
+ PD=5.5e-07 PS=1.52e-06
mXI9.XI166.XI0.XI0.MM2 N_XI9.XI166.XI0.NET12_XI9.XI166.XI0.XI0.MM2_d
+ N_XI9.G13_XI9.XI166.XI0.XI0.MM2_g N_VSS_XI9.XI166.XI0.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.375e-13 AS=2.55e-13
+ PD=5.5e-07 PS=1.52e-06
mXI9.XI165.XI0.XI0.MM2 N_XI9.XI165.XI0.NET12_XI9.XI165.XI0.XI0.MM2_d
+ N_XI9.G12_XI9.XI165.XI0.XI0.MM2_g N_VSS_XI9.XI165.XI0.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.375e-13 AS=2.55e-13
+ PD=5.5e-07 PS=1.52e-06
mXI9.XI159.XI0.XI0.MM2 N_XI9.XI159.XI0.NET12_XI9.XI159.XI0.XI0.MM2_d
+ N_XI9.G11_XI9.XI159.XI0.XI0.MM2_g N_VSS_XI9.XI159.XI0.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.375e-13 AS=2.55e-13
+ PD=5.5e-07 PS=1.52e-06
mXI9.XI160.XI0.XI0.MM2 N_XI9.XI160.XI0.NET12_XI9.XI160.XI0.XI0.MM2_d
+ N_XI9.G10_XI9.XI160.XI0.XI0.MM2_g N_VSS_XI9.XI160.XI0.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.375e-13 AS=2.55e-13
+ PD=5.5e-07 PS=1.52e-06
mXI9.XI161.XI0.XI0.MM2 N_XI9.XI161.XI0.NET12_XI9.XI161.XI0.XI0.MM2_d
+ N_XI9.G9_XI9.XI161.XI0.XI0.MM2_g N_VSS_XI9.XI161.XI0.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.375e-13 AS=2.55e-13
+ PD=5.5e-07 PS=1.52e-06
mXI9.XI162.XI0.XI0.MM2 N_XI9.XI162.XI0.NET12_XI9.XI162.XI0.XI0.MM2_d
+ N_XI9.G8_XI9.XI162.XI0.XI0.MM2_g N_VSS_XI9.XI162.XI0.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.375e-13 AS=2.55e-13
+ PD=5.5e-07 PS=1.52e-06
mXI9.XI121.XI0.XI0.MM2 N_XI9.XI121.XI0.NET12_XI9.XI121.XI0.XI0.MM2_d
+ N_XI9.G7_XI9.XI121.XI0.XI0.MM2_g N_VSS_XI9.XI121.XI0.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.375e-13 AS=2.55e-13
+ PD=5.5e-07 PS=1.52e-06
mXI9.XI120.XI0.XI0.MM2 N_XI9.XI120.XI0.NET12_XI9.XI120.XI0.XI0.MM2_d
+ N_XI9.G6_XI9.XI120.XI0.XI0.MM2_g N_VSS_XI9.XI120.XI0.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.375e-13 AS=2.55e-13
+ PD=5.5e-07 PS=1.52e-06
mXI9.XI119.XI0.XI0.MM2 N_XI9.XI119.XI0.NET12_XI9.XI119.XI0.XI0.MM2_d
+ N_XI9.G5_XI9.XI119.XI0.XI0.MM2_g N_VSS_XI9.XI119.XI0.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.375e-13 AS=2.55e-13
+ PD=5.5e-07 PS=1.52e-06
mXI9.XI118.XI0.XI0.MM2 N_XI9.XI118.XI0.NET12_XI9.XI118.XI0.XI0.MM2_d
+ N_XI9.G4_XI9.XI118.XI0.XI0.MM2_g N_VSS_XI9.XI118.XI0.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.375e-13 AS=2.55e-13
+ PD=5.5e-07 PS=1.52e-06
mXI9.XI91.XI0.XI0.MM2 N_XI9.XI91.XI0.NET12_XI9.XI91.XI0.XI0.MM2_d
+ N_XI9.G3_XI9.XI91.XI0.XI0.MM2_g N_VSS_XI9.XI91.XI0.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.375e-13 AS=2.55e-13
+ PD=5.5e-07 PS=1.52e-06
mXI9.XI90.XI0.XI0.MM2 N_XI9.XI90.XI0.NET12_XI9.XI90.XI0.XI0.MM2_d
+ N_XI9.G2_XI9.XI90.XI0.XI0.MM2_g N_VSS_XI9.XI90.XI0.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.375e-13 AS=2.55e-13
+ PD=5.5e-07 PS=1.52e-06
mXI9.XI89.XI0.XI0.MM2 N_XI9.XI89.XI0.NET12_XI9.XI89.XI0.XI0.MM2_d
+ N_XI9.G1_XI9.XI89.XI0.XI0.MM2_g N_VSS_XI9.XI89.XI0.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.375e-13 AS=2.55e-13
+ PD=5.5e-07 PS=1.52e-06
mXI9.XI168.XI0.XI1.MM2 N_XI9.NET298_XI9.XI168.XI0.XI1.MM2_d
+ N_XI9.XI168.XI0.NET12_XI9.XI168.XI0.XI1.MM2_g N_VSS_XI9.XI168.XI0.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI9.XI167.XI0.XI1.MM2 N_XI9.NET138_XI9.XI167.XI0.XI1.MM2_d
+ N_XI9.XI167.XI0.NET12_XI9.XI167.XI0.XI1.MM2_g N_VSS_XI9.XI167.XI0.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI9.XI166.XI0.XI1.MM2 N_XI9.NET208_XI9.XI166.XI0.XI1.MM2_d
+ N_XI9.XI166.XI0.NET12_XI9.XI166.XI0.XI1.MM2_g N_VSS_XI9.XI166.XI0.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI9.XI165.XI0.XI1.MM2 N_XI9.NET202_XI9.XI165.XI0.XI1.MM2_d
+ N_XI9.XI165.XI0.NET12_XI9.XI165.XI0.XI1.MM2_g N_VSS_XI9.XI165.XI0.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI9.XI159.XI0.XI1.MM2 N_XI9.NET198_XI9.XI159.XI0.XI1.MM2_d
+ N_XI9.XI159.XI0.NET12_XI9.XI159.XI0.XI1.MM2_g N_VSS_XI9.XI159.XI0.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI9.XI160.XI0.XI1.MM2 N_XI9.NET102_XI9.XI160.XI0.XI1.MM2_d
+ N_XI9.XI160.XI0.NET12_XI9.XI160.XI0.XI1.MM2_g N_VSS_XI9.XI160.XI0.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI9.XI161.XI0.XI1.MM2 N_XI9.NET108_XI9.XI161.XI0.XI1.MM2_d
+ N_XI9.XI161.XI0.NET12_XI9.XI161.XI0.XI1.MM2_g N_VSS_XI9.XI161.XI0.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI9.XI162.XI0.XI1.MM2 N_XI9.NET96_XI9.XI162.XI0.XI1.MM2_d
+ N_XI9.XI162.XI0.NET12_XI9.XI162.XI0.XI1.MM2_g N_VSS_XI9.XI162.XI0.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI9.XI121.XI0.XI1.MM2 N_XI9.NET153_XI9.XI121.XI0.XI1.MM2_d
+ N_XI9.XI121.XI0.NET12_XI9.XI121.XI0.XI1.MM2_g N_VSS_XI9.XI121.XI0.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI9.XI120.XI0.XI1.MM2 N_XI9.NET54_XI9.XI120.XI0.XI1.MM2_d
+ N_XI9.XI120.XI0.NET12_XI9.XI120.XI0.XI1.MM2_g N_VSS_XI9.XI120.XI0.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI9.XI119.XI0.XI1.MM2 N_XI9.NET66_XI9.XI119.XI0.XI1.MM2_d
+ N_XI9.XI119.XI0.NET12_XI9.XI119.XI0.XI1.MM2_g N_VSS_XI9.XI119.XI0.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI9.XI118.XI0.XI1.MM2 N_XI9.NET72_XI9.XI118.XI0.XI1.MM2_d
+ N_XI9.XI118.XI0.NET12_XI9.XI118.XI0.XI1.MM2_g N_VSS_XI9.XI118.XI0.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI9.XI91.XI0.XI1.MM2 N_XI9.NET60_XI9.XI91.XI0.XI1.MM2_d
+ N_XI9.XI91.XI0.NET12_XI9.XI91.XI0.XI1.MM2_g N_VSS_XI9.XI91.XI0.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI9.XI90.XI0.XI1.MM2 N_XI9.NET183_XI9.XI90.XI0.XI1.MM2_d
+ N_XI9.XI90.XI0.NET12_XI9.XI90.XI0.XI1.MM2_g N_VSS_XI9.XI90.XI0.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI9.XI89.XI0.XI1.MM2 N_XI9.NET178_XI9.XI89.XI0.XI1.MM2_d
+ N_XI9.XI89.XI0.NET12_XI9.XI89.XI0.XI1.MM2_g N_VSS_XI9.XI89.XI0.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI26.MM2 N_NET218_XI26.MM2_d N_CLK_XI26.MM2_g N_VSS_XI26.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI27.MM2 N_NET214_XI27.MM2_d N_NET218_XI27.MM2_g N_VSS_XI27.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI9.XI182.XI4.MM2 N_XI9.XI182.NET39_XI9.XI182.XI4.MM2_d
+ N_XI9.NET298_XI9.XI182.XI4.MM2_g N_VSS_XI9.XI182.XI4.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI9.XI181.XI4.MM2 N_XI9.XI181.NET39_XI9.XI181.XI4.MM2_d
+ N_XI9.NET138_XI9.XI181.XI4.MM2_g N_VSS_XI9.XI181.XI4.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI9.XI180.XI4.MM2 N_XI9.XI180.NET39_XI9.XI180.XI4.MM2_d
+ N_XI9.NET208_XI9.XI180.XI4.MM2_g N_VSS_XI9.XI180.XI4.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI9.XI179.XI9.MM2 N_XI9.XI179.NET43_XI9.XI179.XI9.MM2_d
+ N_XI9.NET202_XI9.XI179.XI9.MM2_g N_VSS_XI9.XI179.XI9.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI9.XI178.XI4.MM2 N_XI9.XI178.NET39_XI9.XI178.XI4.MM2_d
+ N_XI9.NET198_XI9.XI178.XI4.MM2_g N_VSS_XI9.XI178.XI4.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI9.XI177.XI4.MM2 N_XI9.XI177.NET39_XI9.XI177.XI4.MM2_d
+ N_XI9.NET102_XI9.XI177.XI4.MM2_g N_VSS_XI9.XI177.XI4.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI9.XI176.XI4.MM2 N_XI9.XI176.NET39_XI9.XI176.XI4.MM2_d
+ N_XI9.NET108_XI9.XI176.XI4.MM2_g N_VSS_XI9.XI176.XI4.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI9.XI175.XI4.MM2 N_XI9.XI175.NET39_XI9.XI175.XI4.MM2_d
+ N_XI9.NET96_XI9.XI175.XI4.MM2_g N_VSS_XI9.XI175.XI4.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI9.XI174.XI4.MM2 N_XI9.XI174.NET39_XI9.XI174.XI4.MM2_d
+ N_XI9.NET153_XI9.XI174.XI4.MM2_g N_VSS_XI9.XI174.XI4.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI9.XI173.XI4.MM2 N_XI9.XI173.NET39_XI9.XI173.XI4.MM2_d
+ N_XI9.NET54_XI9.XI173.XI4.MM2_g N_VSS_XI9.XI173.XI4.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI9.XI172.XI4.MM2 N_XI9.XI172.NET39_XI9.XI172.XI4.MM2_d
+ N_XI9.NET66_XI9.XI172.XI4.MM2_g N_VSS_XI9.XI172.XI4.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI9.XI171.XI4.MM2 N_XI9.XI171.NET39_XI9.XI171.XI4.MM2_d
+ N_XI9.NET72_XI9.XI171.XI4.MM2_g N_VSS_XI9.XI171.XI4.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI9.XI170.XI4.MM2 N_XI9.XI170.NET39_XI9.XI170.XI4.MM2_d
+ N_XI9.NET60_XI9.XI170.XI4.MM2_g N_VSS_XI9.XI170.XI4.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI9.XI96.XI4.MM2 N_XI9.XI96.NET39_XI9.XI96.XI4.MM2_d
+ N_XI9.NET183_XI9.XI96.XI4.MM2_g N_VSS_XI9.XI96.XI4.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI9.XI93.XI4.MM2 N_XI9.XI93.NET39_XI9.XI93.XI4.MM2_d
+ N_XI9.NET178_XI9.XI93.XI4.MM2_g N_VSS_XI9.XI93.XI4.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI9.XI182.MM7 N_XI9.XI182.NET10_XI9.XI182.MM7_d
+ N_XI9.XI182.NET39_XI9.XI182.MM7_g N_VSS_XI9.XI182.MM7_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.2375e-13 AS=3.225e-13
+ PD=8.95e-07 PS=1.79e-06
mXI9.XI181.MM7 N_XI9.XI181.NET10_XI9.XI181.MM7_d
+ N_XI9.XI181.NET39_XI9.XI181.MM7_g N_VSS_XI9.XI181.MM7_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.2375e-13 AS=3.225e-13
+ PD=8.95e-07 PS=1.79e-06
mXI9.XI180.MM7 N_XI9.XI180.NET10_XI9.XI180.MM7_d
+ N_XI9.XI180.NET39_XI9.XI180.MM7_g N_VSS_XI9.XI180.MM7_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.2375e-13 AS=3.225e-13
+ PD=8.95e-07 PS=1.79e-06
mXI9.XI179.MM2 N_XI9.XI179.NET10_XI9.XI179.MM2_d
+ N_XI9.XI179.NET43_XI9.XI179.MM2_g N_VSS_XI9.XI179.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.2375e-13 AS=3.225e-13
+ PD=8.95e-07 PS=1.79e-06
mXI9.XI178.MM7 N_XI9.XI178.NET10_XI9.XI178.MM7_d
+ N_XI9.XI178.NET39_XI9.XI178.MM7_g N_VSS_XI9.XI178.MM7_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.2375e-13 AS=3.225e-13
+ PD=8.95e-07 PS=1.79e-06
mXI9.XI177.MM7 N_XI9.XI177.NET10_XI9.XI177.MM7_d
+ N_XI9.XI177.NET39_XI9.XI177.MM7_g N_VSS_XI9.XI177.MM7_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.2375e-13 AS=3.225e-13
+ PD=8.95e-07 PS=1.79e-06
mXI9.XI176.MM7 N_XI9.XI176.NET10_XI9.XI176.MM7_d
+ N_XI9.XI176.NET39_XI9.XI176.MM7_g N_VSS_XI9.XI176.MM7_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.2375e-13 AS=3.225e-13
+ PD=8.95e-07 PS=1.79e-06
mXI9.XI175.MM7 N_XI9.XI175.NET10_XI9.XI175.MM7_d
+ N_XI9.XI175.NET39_XI9.XI175.MM7_g N_VSS_XI9.XI175.MM7_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.2375e-13 AS=3.225e-13
+ PD=8.95e-07 PS=1.79e-06
mXI9.XI174.MM7 N_XI9.XI174.NET10_XI9.XI174.MM7_d
+ N_XI9.XI174.NET39_XI9.XI174.MM7_g N_VSS_XI9.XI174.MM7_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.2375e-13 AS=3.225e-13
+ PD=8.95e-07 PS=1.79e-06
mXI9.XI173.MM7 N_XI9.XI173.NET10_XI9.XI173.MM7_d
+ N_XI9.XI173.NET39_XI9.XI173.MM7_g N_VSS_XI9.XI173.MM7_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.2375e-13 AS=3.225e-13
+ PD=8.95e-07 PS=1.79e-06
mXI9.XI172.MM7 N_XI9.XI172.NET10_XI9.XI172.MM7_d
+ N_XI9.XI172.NET39_XI9.XI172.MM7_g N_VSS_XI9.XI172.MM7_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.2375e-13 AS=3.225e-13
+ PD=8.95e-07 PS=1.79e-06
mXI9.XI171.MM7 N_XI9.XI171.NET10_XI9.XI171.MM7_d
+ N_XI9.XI171.NET39_XI9.XI171.MM7_g N_VSS_XI9.XI171.MM7_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.2375e-13 AS=3.225e-13
+ PD=8.95e-07 PS=1.79e-06
mXI9.XI170.MM7 N_XI9.XI170.NET10_XI9.XI170.MM7_d
+ N_XI9.XI170.NET39_XI9.XI170.MM7_g N_VSS_XI9.XI170.MM7_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.2375e-13 AS=3.225e-13
+ PD=8.95e-07 PS=1.79e-06
mXI9.XI96.MM7 N_XI9.XI96.NET10_XI9.XI96.MM7_d N_XI9.XI96.NET39_XI9.XI96.MM7_g
+ N_VSS_XI9.XI96.MM7_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.2375e-13 AS=3.225e-13 PD=8.95e-07 PS=1.79e-06
mXI9.XI93.MM7 N_XI9.XI93.NET10_XI9.XI93.MM7_d N_XI9.XI93.NET39_XI9.XI93.MM7_g
+ N_VSS_XI9.XI93.MM7_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.2375e-13 AS=3.225e-13 PD=8.95e-07 PS=1.79e-06
mXI9.XI182.MM2 N_NET177_XI9.XI182.MM2_d N_XI9.XI182.NET43_XI9.XI182.MM2_g
+ N_XI9.XI182.NET10_XI9.XI182.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=4.75e-13 AS=2.2375e-13 PD=1.9e-06 PS=8.95e-07
mXI9.XI181.MM2 N_NET178_XI9.XI181.MM2_d N_XI9.XI181.NET43_XI9.XI181.MM2_g
+ N_XI9.XI181.NET10_XI9.XI181.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=4.75e-13 AS=2.2375e-13 PD=1.9e-06 PS=8.95e-07
mXI9.XI180.MM2 N_NET179_XI9.XI180.MM2_d N_XI9.XI180.NET43_XI9.XI180.MM2_g
+ N_XI9.XI180.NET10_XI9.XI180.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=4.75e-13 AS=2.2375e-13 PD=1.9e-06 PS=8.95e-07
mXI9.XI179.MM7 N_NET180_XI9.XI179.MM7_d N_XI9.XI179.NET39_XI9.XI179.MM7_g
+ N_XI9.XI179.NET10_XI9.XI179.MM7_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=4.75e-13 AS=2.2375e-13 PD=1.9e-06 PS=8.95e-07
mXI9.XI178.MM2 N_NET181_XI9.XI178.MM2_d N_XI9.XI178.NET43_XI9.XI178.MM2_g
+ N_XI9.XI178.NET10_XI9.XI178.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=4.75e-13 AS=2.2375e-13 PD=1.9e-06 PS=8.95e-07
mXI9.XI177.MM2 N_NET182_XI9.XI177.MM2_d N_XI9.XI177.NET43_XI9.XI177.MM2_g
+ N_XI9.XI177.NET10_XI9.XI177.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=4.75e-13 AS=2.2375e-13 PD=1.9e-06 PS=8.95e-07
mXI9.XI176.MM2 N_NET183_XI9.XI176.MM2_d N_XI9.XI176.NET43_XI9.XI176.MM2_g
+ N_XI9.XI176.NET10_XI9.XI176.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=4.75e-13 AS=2.2375e-13 PD=1.9e-06 PS=8.95e-07
mXI9.XI175.MM2 N_NET184_XI9.XI175.MM2_d N_XI9.XI175.NET43_XI9.XI175.MM2_g
+ N_XI9.XI175.NET10_XI9.XI175.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=4.75e-13 AS=2.2375e-13 PD=1.9e-06 PS=8.95e-07
mXI9.XI174.MM2 N_NET185_XI9.XI174.MM2_d N_XI9.XI174.NET43_XI9.XI174.MM2_g
+ N_XI9.XI174.NET10_XI9.XI174.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=4.75e-13 AS=2.2375e-13 PD=1.9e-06 PS=8.95e-07
mXI9.XI173.MM2 N_NET186_XI9.XI173.MM2_d N_XI9.XI173.NET43_XI9.XI173.MM2_g
+ N_XI9.XI173.NET10_XI9.XI173.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=4.75e-13 AS=2.2375e-13 PD=1.9e-06 PS=8.95e-07
mXI9.XI172.MM2 N_NET187_XI9.XI172.MM2_d N_XI9.XI172.NET43_XI9.XI172.MM2_g
+ N_XI9.XI172.NET10_XI9.XI172.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=4.75e-13 AS=2.2375e-13 PD=1.9e-06 PS=8.95e-07
mXI9.XI171.MM2 N_NET188_XI9.XI171.MM2_d N_XI9.XI171.NET43_XI9.XI171.MM2_g
+ N_XI9.XI171.NET10_XI9.XI171.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=4.75e-13 AS=2.2375e-13 PD=1.9e-06 PS=8.95e-07
mXI9.XI170.MM2 N_NET189_XI9.XI170.MM2_d N_XI9.XI170.NET43_XI9.XI170.MM2_g
+ N_XI9.XI170.NET10_XI9.XI170.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=4.75e-13 AS=2.2375e-13 PD=1.9e-06 PS=8.95e-07
mXI9.XI96.MM2 N_NET190_XI9.XI96.MM2_d N_XI9.XI96.NET43_XI9.XI96.MM2_g
+ N_XI9.XI96.NET10_XI9.XI96.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=4.75e-13 AS=2.2375e-13 PD=1.9e-06 PS=8.95e-07
mXI9.XI93.MM2 N_NET191_XI9.XI93.MM2_d N_XI9.XI93.NET43_XI9.XI93.MM2_g
+ N_XI9.XI93.NET10_XI9.XI93.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=4.75e-13 AS=2.2375e-13 PD=1.9e-06 PS=8.95e-07
mXI28.MM2 N_NET210_XI28.MM2_d N_NET214_XI28.MM2_g N_VSS_XI28.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=3e-06 AD=1.47e-12 AS=1.47e-12
+ PD=3.98e-06 PS=3.98e-06
mXI29.MM2 N_NET222_XI29.MM2_d N_NET210_XI29.MM2_g N_VSS_XI29.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=3e-06 AD=1.47e-12 AS=1.47e-12
+ PD=3.98e-06 PS=3.98e-06
mXI9.XI182.MM0 N_NET177_XI9.XI182.MM0_d N_XI9.P16_XI9.XI182.MM0_g
+ N_XI9.XI182.NET6_XI9.XI182.MM0_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=4.75e-13 AS=1.8125e-13 PD=1.9e-06 PS=7.25e-07
mXI9.XI181.MM0 N_NET178_XI9.XI181.MM0_d N_XI9.P15_XI9.XI181.MM0_g
+ N_XI9.XI181.NET6_XI9.XI181.MM0_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=4.75e-13 AS=1.8125e-13 PD=1.9e-06 PS=7.25e-07
mXI9.XI180.MM0 N_NET179_XI9.XI180.MM0_d N_XI9.P14_XI9.XI180.MM0_g
+ N_XI9.XI180.NET6_XI9.XI180.MM0_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=4.75e-13 AS=1.8125e-13 PD=1.9e-06 PS=7.25e-07
mXI9.XI179.MM6 N_NET180_XI9.XI179.MM6_d N_XI9.P13_XI9.XI179.MM6_g
+ N_XI9.XI179.NET6_XI9.XI179.MM6_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=4.75e-13 AS=1.8125e-13 PD=1.9e-06 PS=7.25e-07
mXI9.XI178.MM0 N_NET181_XI9.XI178.MM0_d N_XI9.P12_XI9.XI178.MM0_g
+ N_XI9.XI178.NET6_XI9.XI178.MM0_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=4.75e-13 AS=1.8125e-13 PD=1.9e-06 PS=7.25e-07
mXI9.XI177.MM0 N_NET182_XI9.XI177.MM0_d N_XI9.P11_XI9.XI177.MM0_g
+ N_XI9.XI177.NET6_XI9.XI177.MM0_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=4.75e-13 AS=1.8125e-13 PD=1.9e-06 PS=7.25e-07
mXI9.XI176.MM0 N_NET183_XI9.XI176.MM0_d N_XI9.P10_XI9.XI176.MM0_g
+ N_XI9.XI176.NET6_XI9.XI176.MM0_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=4.75e-13 AS=1.8125e-13 PD=1.9e-06 PS=7.25e-07
mXI9.XI175.MM0 N_NET184_XI9.XI175.MM0_d N_XI9.P9_XI9.XI175.MM0_g
+ N_XI9.XI175.NET6_XI9.XI175.MM0_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=4.75e-13 AS=1.8125e-13 PD=1.9e-06 PS=7.25e-07
mXI9.XI174.MM0 N_NET185_XI9.XI174.MM0_d N_XI9.P8_XI9.XI174.MM0_g
+ N_XI9.XI174.NET6_XI9.XI174.MM0_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=4.75e-13 AS=1.8125e-13 PD=1.9e-06 PS=7.25e-07
mXI9.XI173.MM0 N_NET186_XI9.XI173.MM0_d N_XI9.P7_XI9.XI173.MM0_g
+ N_XI9.XI173.NET6_XI9.XI173.MM0_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=4.75e-13 AS=1.8125e-13 PD=1.9e-06 PS=7.25e-07
mXI9.XI172.MM0 N_NET187_XI9.XI172.MM0_d N_XI9.P6_XI9.XI172.MM0_g
+ N_XI9.XI172.NET6_XI9.XI172.MM0_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=4.75e-13 AS=1.8125e-13 PD=1.9e-06 PS=7.25e-07
mXI9.XI171.MM0 N_NET188_XI9.XI171.MM0_d N_XI9.P5_XI9.XI171.MM0_g
+ N_XI9.XI171.NET6_XI9.XI171.MM0_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=4.75e-13 AS=1.8125e-13 PD=1.9e-06 PS=7.25e-07
mXI9.XI170.MM0 N_NET189_XI9.XI170.MM0_d N_XI9.P4_XI9.XI170.MM0_g
+ N_XI9.XI170.NET6_XI9.XI170.MM0_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=4.75e-13 AS=1.8125e-13 PD=1.9e-06 PS=7.25e-07
mXI9.XI96.MM0 N_NET190_XI9.XI96.MM0_d N_XI9.P3_XI9.XI96.MM0_g
+ N_XI9.XI96.NET6_XI9.XI96.MM0_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=4.75e-13 AS=1.8125e-13 PD=1.9e-06 PS=7.25e-07
mXI9.XI93.MM0 N_NET191_XI9.XI93.MM0_d N_XI9.P2_XI9.XI93.MM0_g
+ N_XI9.XI93.NET6_XI9.XI93.MM0_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=4.75e-13 AS=1.8125e-13 PD=1.9e-06 PS=7.25e-07
mXI9.XI182.MM6 N_XI9.XI182.NET6_XI9.XI182.MM6_d N_XI9.NET298_XI9.XI182.MM6_g
+ N_VSS_XI9.XI182.MM6_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=1.8125e-13 AS=2.575e-13 PD=7.25e-07 PS=1.53e-06
mXI9.XI181.MM6 N_XI9.XI181.NET6_XI9.XI181.MM6_d N_XI9.NET138_XI9.XI181.MM6_g
+ N_VSS_XI9.XI181.MM6_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=1.8125e-13 AS=2.575e-13 PD=7.25e-07 PS=1.53e-06
mXI9.XI180.MM6 N_XI9.XI180.NET6_XI9.XI180.MM6_d N_XI9.NET208_XI9.XI180.MM6_g
+ N_VSS_XI9.XI180.MM6_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=1.8125e-13 AS=2.575e-13 PD=7.25e-07 PS=1.53e-06
mXI9.XI179.MM0 N_XI9.XI179.NET6_XI9.XI179.MM0_d N_XI9.NET202_XI9.XI179.MM0_g
+ N_VSS_XI9.XI179.MM0_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=1.8125e-13 AS=2.575e-13 PD=7.25e-07 PS=1.53e-06
mXI9.XI178.MM6 N_XI9.XI178.NET6_XI9.XI178.MM6_d N_XI9.NET198_XI9.XI178.MM6_g
+ N_VSS_XI9.XI178.MM6_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=1.8125e-13 AS=2.575e-13 PD=7.25e-07 PS=1.53e-06
mXI9.XI177.MM6 N_XI9.XI177.NET6_XI9.XI177.MM6_d N_XI9.NET102_XI9.XI177.MM6_g
+ N_VSS_XI9.XI177.MM6_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=1.8125e-13 AS=2.575e-13 PD=7.25e-07 PS=1.53e-06
mXI9.XI176.MM6 N_XI9.XI176.NET6_XI9.XI176.MM6_d N_XI9.NET108_XI9.XI176.MM6_g
+ N_VSS_XI9.XI176.MM6_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=1.8125e-13 AS=2.575e-13 PD=7.25e-07 PS=1.53e-06
mXI9.XI175.MM6 N_XI9.XI175.NET6_XI9.XI175.MM6_d N_XI9.NET96_XI9.XI175.MM6_g
+ N_VSS_XI9.XI175.MM6_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=1.8125e-13 AS=2.575e-13 PD=7.25e-07 PS=1.53e-06
mXI9.XI174.MM6 N_XI9.XI174.NET6_XI9.XI174.MM6_d N_XI9.NET153_XI9.XI174.MM6_g
+ N_VSS_XI9.XI174.MM6_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=1.8125e-13 AS=2.575e-13 PD=7.25e-07 PS=1.53e-06
mXI9.XI173.MM6 N_XI9.XI173.NET6_XI9.XI173.MM6_d N_XI9.NET54_XI9.XI173.MM6_g
+ N_VSS_XI9.XI173.MM6_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=1.8125e-13 AS=2.575e-13 PD=7.25e-07 PS=1.53e-06
mXI9.XI172.MM6 N_XI9.XI172.NET6_XI9.XI172.MM6_d N_XI9.NET66_XI9.XI172.MM6_g
+ N_VSS_XI9.XI172.MM6_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=1.8125e-13 AS=2.575e-13 PD=7.25e-07 PS=1.53e-06
mXI9.XI171.MM6 N_XI9.XI171.NET6_XI9.XI171.MM6_d N_XI9.NET72_XI9.XI171.MM6_g
+ N_VSS_XI9.XI171.MM6_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=1.8125e-13 AS=2.575e-13 PD=7.25e-07 PS=1.53e-06
mXI9.XI170.MM6 N_XI9.XI170.NET6_XI9.XI170.MM6_d N_XI9.NET60_XI9.XI170.MM6_g
+ N_VSS_XI9.XI170.MM6_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=1.8125e-13 AS=2.575e-13 PD=7.25e-07 PS=1.53e-06
mXI9.XI96.MM6 N_XI9.XI96.NET6_XI9.XI96.MM6_d N_XI9.NET183_XI9.XI96.MM6_g
+ N_VSS_XI9.XI96.MM6_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=1.8125e-13 AS=2.575e-13 PD=7.25e-07 PS=1.53e-06
mXI9.XI93.MM6 N_XI9.XI93.NET6_XI9.XI93.MM6_d N_XI9.NET178_XI9.XI93.MM6_g
+ N_VSS_XI9.XI93.MM6_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=1.8125e-13 AS=2.575e-13 PD=7.25e-07 PS=1.53e-06
mXI9.XI182.XI9.MM2 N_XI9.XI182.NET43_XI9.XI182.XI9.MM2_d
+ N_XI9.P16_XI9.XI182.XI9.MM2_g N_VSS_XI9.XI182.XI9.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI9.XI181.XI9.MM2 N_XI9.XI181.NET43_XI9.XI181.XI9.MM2_d
+ N_XI9.P15_XI9.XI181.XI9.MM2_g N_VSS_XI9.XI181.XI9.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI9.XI180.XI9.MM2 N_XI9.XI180.NET43_XI9.XI180.XI9.MM2_d
+ N_XI9.P14_XI9.XI180.XI9.MM2_g N_VSS_XI9.XI180.XI9.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI9.XI179.XI4.MM2 N_XI9.XI179.NET39_XI9.XI179.XI4.MM2_d
+ N_XI9.P13_XI9.XI179.XI4.MM2_g N_VSS_XI9.XI179.XI4.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI9.XI178.XI9.MM2 N_XI9.XI178.NET43_XI9.XI178.XI9.MM2_d
+ N_XI9.P12_XI9.XI178.XI9.MM2_g N_VSS_XI9.XI178.XI9.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI9.XI177.XI9.MM2 N_XI9.XI177.NET43_XI9.XI177.XI9.MM2_d
+ N_XI9.P11_XI9.XI177.XI9.MM2_g N_VSS_XI9.XI177.XI9.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI9.XI176.XI9.MM2 N_XI9.XI176.NET43_XI9.XI176.XI9.MM2_d
+ N_XI9.P10_XI9.XI176.XI9.MM2_g N_VSS_XI9.XI176.XI9.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI9.XI175.XI9.MM2 N_XI9.XI175.NET43_XI9.XI175.XI9.MM2_d
+ N_XI9.P9_XI9.XI175.XI9.MM2_g N_VSS_XI9.XI175.XI9.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI9.XI174.XI9.MM2 N_XI9.XI174.NET43_XI9.XI174.XI9.MM2_d
+ N_XI9.P8_XI9.XI174.XI9.MM2_g N_VSS_XI9.XI174.XI9.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI9.XI173.XI9.MM2 N_XI9.XI173.NET43_XI9.XI173.XI9.MM2_d
+ N_XI9.P7_XI9.XI173.XI9.MM2_g N_VSS_XI9.XI173.XI9.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI9.XI172.XI9.MM2 N_XI9.XI172.NET43_XI9.XI172.XI9.MM2_d
+ N_XI9.P6_XI9.XI172.XI9.MM2_g N_VSS_XI9.XI172.XI9.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI9.XI171.XI9.MM2 N_XI9.XI171.NET43_XI9.XI171.XI9.MM2_d
+ N_XI9.P5_XI9.XI171.XI9.MM2_g N_VSS_XI9.XI171.XI9.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI9.XI170.XI9.MM2 N_XI9.XI170.NET43_XI9.XI170.XI9.MM2_d
+ N_XI9.P4_XI9.XI170.XI9.MM2_g N_VSS_XI9.XI170.XI9.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI9.XI96.XI9.MM2 N_XI9.XI96.NET43_XI9.XI96.XI9.MM2_d
+ N_XI9.P3_XI9.XI96.XI9.MM2_g N_VSS_XI9.XI96.XI9.MM2_s N_VSS_XI10.XI0.XI0.MM2_b
+ N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI9.XI93.XI9.MM2 N_XI9.XI93.NET43_XI9.XI93.XI9.MM2_d
+ N_XI9.P2_XI9.XI93.XI9.MM2_g N_VSS_XI9.XI93.XI9.MM2_s N_VSS_XI10.XI0.XI0.MM2_b
+ N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI16.XI30.XI1.MM0 N_XI16.XI30.XI1.NET036_XI16.XI30.XI1.MM0_d
+ N_NET198_XI16.XI30.XI1.MM0_g N_VSS_XI16.XI30.XI1.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.375e-13 AS=2.45e-13
+ PD=5.5e-07 PS=1.48e-06
mXI16.XI29.XI1.MM0 N_XI16.XI29.XI1.NET036_XI16.XI29.XI1.MM0_d
+ N_NET198_XI16.XI29.XI1.MM0_g N_VSS_XI16.XI29.XI1.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.375e-13 AS=2.45e-13
+ PD=5.5e-07 PS=1.48e-06
mXI16.XI28.XI1.MM0 N_XI16.XI28.XI1.NET036_XI16.XI28.XI1.MM0_d
+ N_NET198_XI16.XI28.XI1.MM0_g N_VSS_XI16.XI28.XI1.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.375e-13 AS=2.45e-13
+ PD=5.5e-07 PS=1.48e-06
mXI16.XI27.XI1.MM0 N_XI16.XI27.XI1.NET036_XI16.XI27.XI1.MM0_d
+ N_NET198_XI16.XI27.XI1.MM0_g N_VSS_XI16.XI27.XI1.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.375e-13 AS=2.45e-13
+ PD=5.5e-07 PS=1.48e-06
mXI16.XI26.XI1.MM0 N_XI16.XI26.XI1.NET036_XI16.XI26.XI1.MM0_d
+ N_NET198_XI16.XI26.XI1.MM0_g N_VSS_XI16.XI26.XI1.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.375e-13 AS=2.45e-13
+ PD=5.5e-07 PS=1.48e-06
mXI16.XI25.XI1.MM0 N_XI16.XI25.XI1.NET036_XI16.XI25.XI1.MM0_d
+ N_NET198_XI16.XI25.XI1.MM0_g N_VSS_XI16.XI25.XI1.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.375e-13 AS=2.45e-13
+ PD=5.5e-07 PS=1.48e-06
mXI16.XI24.XI1.MM0 N_XI16.XI24.XI1.NET036_XI16.XI24.XI1.MM0_d
+ N_NET198_XI16.XI24.XI1.MM0_g N_VSS_XI16.XI24.XI1.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.375e-13 AS=2.45e-13
+ PD=5.5e-07 PS=1.48e-06
mXI16.XI23.XI1.MM0 N_XI16.XI23.XI1.NET036_XI16.XI23.XI1.MM0_d
+ N_NET198_XI16.XI23.XI1.MM0_g N_VSS_XI16.XI23.XI1.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.375e-13 AS=2.45e-13
+ PD=5.5e-07 PS=1.48e-06
mXI16.XI22.XI1.MM0 N_XI16.XI22.XI1.NET036_XI16.XI22.XI1.MM0_d
+ N_NET198_XI16.XI22.XI1.MM0_g N_VSS_XI16.XI22.XI1.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.375e-13 AS=2.45e-13
+ PD=5.5e-07 PS=1.48e-06
mXI16.XI21.XI1.MM0 N_XI16.XI21.XI1.NET036_XI16.XI21.XI1.MM0_d
+ N_NET198_XI16.XI21.XI1.MM0_g N_VSS_XI16.XI21.XI1.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.375e-13 AS=2.45e-13
+ PD=5.5e-07 PS=1.48e-06
mXI16.XI20.XI1.MM0 N_XI16.XI20.XI1.NET036_XI16.XI20.XI1.MM0_d
+ N_NET198_XI16.XI20.XI1.MM0_g N_VSS_XI16.XI20.XI1.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.375e-13 AS=2.45e-13
+ PD=5.5e-07 PS=1.48e-06
mXI16.XI19.XI1.MM0 N_XI16.XI19.XI1.NET036_XI16.XI19.XI1.MM0_d
+ N_NET198_XI16.XI19.XI1.MM0_g N_VSS_XI16.XI19.XI1.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.375e-13 AS=2.45e-13
+ PD=5.5e-07 PS=1.48e-06
mXI16.XI18.XI1.MM0 N_XI16.XI18.XI1.NET036_XI16.XI18.XI1.MM0_d
+ N_NET198_XI16.XI18.XI1.MM0_g N_VSS_XI16.XI18.XI1.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.375e-13 AS=2.45e-13
+ PD=5.5e-07 PS=1.48e-06
mXI16.XI17.XI1.MM0 N_XI16.XI17.XI1.NET036_XI16.XI17.XI1.MM0_d
+ N_NET198_XI16.XI17.XI1.MM0_g N_VSS_XI16.XI17.XI1.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.375e-13 AS=2.45e-13
+ PD=5.5e-07 PS=1.48e-06
mXI16.XI16.XI1.MM0 N_XI16.XI16.XI1.NET036_XI16.XI16.XI1.MM0_d
+ N_NET198_XI16.XI16.XI1.MM0_g N_VSS_XI16.XI16.XI1.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.375e-13 AS=2.45e-13
+ PD=5.5e-07 PS=1.48e-06
mXI16.XI0.XI1.MM2 N_XI16.XI0.XI1.NET036_XI16.XI0.XI1.MM2_d
+ N_NET198_XI16.XI0.XI1.MM2_g N_VSS_XI16.XI0.XI1.MM2_s N_VSS_XI10.XI0.XI0.MM2_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.375e-13 AS=2.45e-13 PD=5.5e-07 PS=1.48e-06
mXI16.XI30.XI1.MM2 N_XI16.XI30.NET6_XI16.XI30.XI1.MM2_d
+ N_NET177_XI16.XI30.XI1.MM2_g N_XI16.XI30.XI1.NET036_XI16.XI30.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=1.375e-13
+ PD=1.52e-06 PS=5.5e-07
mXI16.XI29.XI1.MM2 N_XI16.XI29.NET6_XI16.XI29.XI1.MM2_d
+ N_NET178_XI16.XI29.XI1.MM2_g N_XI16.XI29.XI1.NET036_XI16.XI29.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=1.375e-13
+ PD=1.52e-06 PS=5.5e-07
mXI16.XI28.XI1.MM2 N_XI16.XI28.NET6_XI16.XI28.XI1.MM2_d
+ N_NET179_XI16.XI28.XI1.MM2_g N_XI16.XI28.XI1.NET036_XI16.XI28.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=1.375e-13
+ PD=1.52e-06 PS=5.5e-07
mXI16.XI27.XI1.MM2 N_XI16.XI27.NET6_XI16.XI27.XI1.MM2_d
+ N_NET180_XI16.XI27.XI1.MM2_g N_XI16.XI27.XI1.NET036_XI16.XI27.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=1.375e-13
+ PD=1.52e-06 PS=5.5e-07
mXI16.XI26.XI1.MM2 N_XI16.XI26.NET6_XI16.XI26.XI1.MM2_d
+ N_NET181_XI16.XI26.XI1.MM2_g N_XI16.XI26.XI1.NET036_XI16.XI26.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=1.375e-13
+ PD=1.52e-06 PS=5.5e-07
mXI16.XI25.XI1.MM2 N_XI16.XI25.NET6_XI16.XI25.XI1.MM2_d
+ N_NET182_XI16.XI25.XI1.MM2_g N_XI16.XI25.XI1.NET036_XI16.XI25.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=1.375e-13
+ PD=1.52e-06 PS=5.5e-07
mXI16.XI24.XI1.MM2 N_XI16.XI24.NET6_XI16.XI24.XI1.MM2_d
+ N_NET183_XI16.XI24.XI1.MM2_g N_XI16.XI24.XI1.NET036_XI16.XI24.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=1.375e-13
+ PD=1.52e-06 PS=5.5e-07
mXI16.XI23.XI1.MM2 N_XI16.XI23.NET6_XI16.XI23.XI1.MM2_d
+ N_NET184_XI16.XI23.XI1.MM2_g N_XI16.XI23.XI1.NET036_XI16.XI23.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=1.375e-13
+ PD=1.52e-06 PS=5.5e-07
mXI16.XI22.XI1.MM2 N_XI16.XI22.NET6_XI16.XI22.XI1.MM2_d
+ N_NET185_XI16.XI22.XI1.MM2_g N_XI16.XI22.XI1.NET036_XI16.XI22.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=1.375e-13
+ PD=1.52e-06 PS=5.5e-07
mXI16.XI21.XI1.MM2 N_XI16.XI21.NET6_XI16.XI21.XI1.MM2_d
+ N_NET186_XI16.XI21.XI1.MM2_g N_XI16.XI21.XI1.NET036_XI16.XI21.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=1.375e-13
+ PD=1.52e-06 PS=5.5e-07
mXI16.XI20.XI1.MM2 N_XI16.XI20.NET6_XI16.XI20.XI1.MM2_d
+ N_NET187_XI16.XI20.XI1.MM2_g N_XI16.XI20.XI1.NET036_XI16.XI20.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=1.375e-13
+ PD=1.52e-06 PS=5.5e-07
mXI16.XI19.XI1.MM2 N_XI16.XI19.NET6_XI16.XI19.XI1.MM2_d
+ N_NET188_XI16.XI19.XI1.MM2_g N_XI16.XI19.XI1.NET036_XI16.XI19.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=1.375e-13
+ PD=1.52e-06 PS=5.5e-07
mXI16.XI18.XI1.MM2 N_XI16.XI18.NET6_XI16.XI18.XI1.MM2_d
+ N_NET189_XI16.XI18.XI1.MM2_g N_XI16.XI18.XI1.NET036_XI16.XI18.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=1.375e-13
+ PD=1.52e-06 PS=5.5e-07
mXI16.XI17.XI1.MM2 N_XI16.XI17.NET6_XI16.XI17.XI1.MM2_d
+ N_NET190_XI16.XI17.XI1.MM2_g N_XI16.XI17.XI1.NET036_XI16.XI17.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=1.375e-13
+ PD=1.52e-06 PS=5.5e-07
mXI16.XI16.XI1.MM2 N_XI16.XI16.NET6_XI16.XI16.XI1.MM2_d
+ N_NET191_XI16.XI16.XI1.MM2_g N_XI16.XI16.XI1.NET036_XI16.XI16.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=1.375e-13
+ PD=1.52e-06 PS=5.5e-07
mXI16.XI0.XI1.MM0 N_XI16.XI0.NET6_XI16.XI0.XI1.MM0_d N_NET192_XI16.XI0.XI1.MM0_g
+ N_XI16.XI0.XI1.NET036_XI16.XI0.XI1.MM0_s N_VSS_XI10.XI0.XI0.MM2_b N_18
+ L=1.8e-07 W=5e-07 AD=2.55e-13 AS=1.375e-13 PD=1.52e-06 PS=5.5e-07
mXI16.XI30.XI0.MM2 N_NET452_XI16.XI30.XI0.MM2_d
+ N_XI16.XI30.NET6_XI16.XI30.XI0.MM2_g N_VSS_XI16.XI30.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI16.XI29.XI0.MM2 N_NET453_XI16.XI29.XI0.MM2_d
+ N_XI16.XI29.NET6_XI16.XI29.XI0.MM2_g N_VSS_XI16.XI29.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI16.XI28.XI0.MM2 N_NET454_XI16.XI28.XI0.MM2_d
+ N_XI16.XI28.NET6_XI16.XI28.XI0.MM2_g N_VSS_XI16.XI28.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI16.XI27.XI0.MM2 N_NET455_XI16.XI27.XI0.MM2_d
+ N_XI16.XI27.NET6_XI16.XI27.XI0.MM2_g N_VSS_XI16.XI27.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI16.XI26.XI0.MM2 N_NET456_XI16.XI26.XI0.MM2_d
+ N_XI16.XI26.NET6_XI16.XI26.XI0.MM2_g N_VSS_XI16.XI26.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI16.XI25.XI0.MM2 N_NET457_XI16.XI25.XI0.MM2_d
+ N_XI16.XI25.NET6_XI16.XI25.XI0.MM2_g N_VSS_XI16.XI25.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI16.XI24.XI0.MM2 N_NET458_XI16.XI24.XI0.MM2_d
+ N_XI16.XI24.NET6_XI16.XI24.XI0.MM2_g N_VSS_XI16.XI24.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI16.XI23.XI0.MM2 N_NET459_XI16.XI23.XI0.MM2_d
+ N_XI16.XI23.NET6_XI16.XI23.XI0.MM2_g N_VSS_XI16.XI23.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI16.XI22.XI0.MM2 N_NET460_XI16.XI22.XI0.MM2_d
+ N_XI16.XI22.NET6_XI16.XI22.XI0.MM2_g N_VSS_XI16.XI22.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI16.XI21.XI0.MM2 N_NET461_XI16.XI21.XI0.MM2_d
+ N_XI16.XI21.NET6_XI16.XI21.XI0.MM2_g N_VSS_XI16.XI21.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI16.XI20.XI0.MM2 N_NET462_XI16.XI20.XI0.MM2_d
+ N_XI16.XI20.NET6_XI16.XI20.XI0.MM2_g N_VSS_XI16.XI20.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI16.XI19.XI0.MM2 N_NET463_XI16.XI19.XI0.MM2_d
+ N_XI16.XI19.NET6_XI16.XI19.XI0.MM2_g N_VSS_XI16.XI19.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI16.XI18.XI0.MM2 N_NET464_XI16.XI18.XI0.MM2_d
+ N_XI16.XI18.NET6_XI16.XI18.XI0.MM2_g N_VSS_XI16.XI18.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI16.XI17.XI0.MM2 N_NET465_XI16.XI17.XI0.MM2_d
+ N_XI16.XI17.NET6_XI16.XI17.XI0.MM2_g N_VSS_XI16.XI17.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI16.XI16.XI0.MM2 N_NET466_XI16.XI16.XI0.MM2_d
+ N_XI16.XI16.NET6_XI16.XI16.XI0.MM2_g N_VSS_XI16.XI16.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI16.XI0.XI0.MM2 N_NET467_XI16.XI0.XI0.MM2_d N_XI16.XI0.NET6_XI16.XI0.XI0.MM2_g
+ N_VSS_XI16.XI0.XI0.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI11.XI30.XI0.MM2 N_XI11.XI30.NET0180_XI11.XI30.XI0.MM2_d
+ N_NET222_XI11.XI30.XI0.MM2_g N_VSS_XI11.XI30.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI29.XI0.MM2 N_XI11.XI29.NET0180_XI11.XI29.XI0.MM2_d
+ N_NET222_XI11.XI29.XI0.MM2_g N_VSS_XI11.XI29.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI31.XI0.MM2 N_XI11.XI31.NET0180_XI11.XI31.XI0.MM2_d
+ N_NET222_XI11.XI31.XI0.MM2_g N_VSS_XI11.XI31.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI28.XI0.MM2 N_XI11.XI28.NET0180_XI11.XI28.XI0.MM2_d
+ N_NET222_XI11.XI28.XI0.MM2_g N_VSS_XI11.XI28.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI25.XI0.MM2 N_XI11.XI25.NET0180_XI11.XI25.XI0.MM2_d
+ N_NET222_XI11.XI25.XI0.MM2_g N_VSS_XI11.XI25.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI26.XI0.MM2 N_XI11.XI26.NET0180_XI11.XI26.XI0.MM2_d
+ N_NET222_XI11.XI26.XI0.MM2_g N_VSS_XI11.XI26.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI24.XI0.MM2 N_XI11.XI24.NET0180_XI11.XI24.XI0.MM2_d
+ N_NET222_XI11.XI24.XI0.MM2_g N_VSS_XI11.XI24.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI27.XI0.MM2 N_XI11.XI27.NET0180_XI11.XI27.XI0.MM2_d
+ N_NET222_XI11.XI27.XI0.MM2_g N_VSS_XI11.XI27.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI22.XI0.MM2 N_XI11.XI22.NET0180_XI11.XI22.XI0.MM2_d
+ N_NET222_XI11.XI22.XI0.MM2_g N_VSS_XI11.XI22.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI21.XI0.MM2 N_XI11.XI21.NET0180_XI11.XI21.XI0.MM2_d
+ N_NET222_XI11.XI21.XI0.MM2_g N_VSS_XI11.XI21.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI23.XI0.MM2 N_XI11.XI23.NET0180_XI11.XI23.XI0.MM2_d
+ N_NET222_XI11.XI23.XI0.MM2_g N_VSS_XI11.XI23.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI19.XI0.MM2 N_XI11.XI19.NET0180_XI11.XI19.XI0.MM2_d
+ N_NET222_XI11.XI19.XI0.MM2_g N_VSS_XI11.XI19.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI20.XI0.MM2 N_XI11.XI20.NET0180_XI11.XI20.XI0.MM2_d
+ N_NET222_XI11.XI20.XI0.MM2_g N_VSS_XI11.XI20.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI18.XI0.MM2 N_XI11.XI18.NET0180_XI11.XI18.XI0.MM2_d
+ N_NET222_XI11.XI18.XI0.MM2_g N_VSS_XI11.XI18.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI17.XI0.MM2 N_XI11.XI17.NET0180_XI11.XI17.XI0.MM2_d
+ N_NET222_XI11.XI17.XI0.MM2_g N_VSS_XI11.XI17.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI0.XI0.MM2 N_XI11.XI0.NET0180_XI11.XI0.XI0.MM2_d
+ N_NET222_XI11.XI0.XI0.MM2_g N_VSS_XI11.XI0.XI0.MM2_s N_VSS_XI10.XI0.XI0.MM2_b
+ N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI11.XI30.XI1.MM2 N_XI11.XI30.NET35_XI11.XI30.XI1.MM2_d
+ N_XI11.XI30.NET0180_XI11.XI30.XI1.MM2_g N_VSS_XI11.XI30.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI29.XI1.MM2 N_XI11.XI29.NET35_XI11.XI29.XI1.MM2_d
+ N_XI11.XI29.NET0180_XI11.XI29.XI1.MM2_g N_VSS_XI11.XI29.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI31.XI1.MM2 N_XI11.XI31.NET35_XI11.XI31.XI1.MM2_d
+ N_XI11.XI31.NET0180_XI11.XI31.XI1.MM2_g N_VSS_XI11.XI31.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI28.XI1.MM2 N_XI11.XI28.NET35_XI11.XI28.XI1.MM2_d
+ N_XI11.XI28.NET0180_XI11.XI28.XI1.MM2_g N_VSS_XI11.XI28.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI25.XI1.MM2 N_XI11.XI25.NET35_XI11.XI25.XI1.MM2_d
+ N_XI11.XI25.NET0180_XI11.XI25.XI1.MM2_g N_VSS_XI11.XI25.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI26.XI1.MM2 N_XI11.XI26.NET35_XI11.XI26.XI1.MM2_d
+ N_XI11.XI26.NET0180_XI11.XI26.XI1.MM2_g N_VSS_XI11.XI26.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI24.XI1.MM2 N_XI11.XI24.NET35_XI11.XI24.XI1.MM2_d
+ N_XI11.XI24.NET0180_XI11.XI24.XI1.MM2_g N_VSS_XI11.XI24.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI27.XI1.MM2 N_XI11.XI27.NET35_XI11.XI27.XI1.MM2_d
+ N_XI11.XI27.NET0180_XI11.XI27.XI1.MM2_g N_VSS_XI11.XI27.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI22.XI1.MM2 N_XI11.XI22.NET35_XI11.XI22.XI1.MM2_d
+ N_XI11.XI22.NET0180_XI11.XI22.XI1.MM2_g N_VSS_XI11.XI22.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI21.XI1.MM2 N_XI11.XI21.NET35_XI11.XI21.XI1.MM2_d
+ N_XI11.XI21.NET0180_XI11.XI21.XI1.MM2_g N_VSS_XI11.XI21.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI23.XI1.MM2 N_XI11.XI23.NET35_XI11.XI23.XI1.MM2_d
+ N_XI11.XI23.NET0180_XI11.XI23.XI1.MM2_g N_VSS_XI11.XI23.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI19.XI1.MM2 N_XI11.XI19.NET35_XI11.XI19.XI1.MM2_d
+ N_XI11.XI19.NET0180_XI11.XI19.XI1.MM2_g N_VSS_XI11.XI19.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI20.XI1.MM2 N_XI11.XI20.NET35_XI11.XI20.XI1.MM2_d
+ N_XI11.XI20.NET0180_XI11.XI20.XI1.MM2_g N_VSS_XI11.XI20.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI18.XI1.MM2 N_XI11.XI18.NET35_XI11.XI18.XI1.MM2_d
+ N_XI11.XI18.NET0180_XI11.XI18.XI1.MM2_g N_VSS_XI11.XI18.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI17.XI1.MM2 N_XI11.XI17.NET35_XI11.XI17.XI1.MM2_d
+ N_XI11.XI17.NET0180_XI11.XI17.XI1.MM2_g N_VSS_XI11.XI17.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI0.XI1.MM2 N_XI11.XI0.NET35_XI11.XI0.XI1.MM2_d
+ N_XI11.XI0.NET0180_XI11.XI0.XI1.MM2_g N_VSS_XI11.XI0.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI30.MM26 N_XI11.XI30.CLKB_XI11.XI30.MM26_d
+ N_XI11.XI30.NET35_XI11.XI30.MM26_g N_VSS_XI11.XI30.MM26_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI29.MM26 N_XI11.XI29.CLKB_XI11.XI29.MM26_d
+ N_XI11.XI29.NET35_XI11.XI29.MM26_g N_VSS_XI11.XI29.MM26_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI31.MM26 N_XI11.XI31.CLKB_XI11.XI31.MM26_d
+ N_XI11.XI31.NET35_XI11.XI31.MM26_g N_VSS_XI11.XI31.MM26_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI28.MM26 N_XI11.XI28.CLKB_XI11.XI28.MM26_d
+ N_XI11.XI28.NET35_XI11.XI28.MM26_g N_VSS_XI11.XI28.MM26_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI25.MM26 N_XI11.XI25.CLKB_XI11.XI25.MM26_d
+ N_XI11.XI25.NET35_XI11.XI25.MM26_g N_VSS_XI11.XI25.MM26_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI26.MM26 N_XI11.XI26.CLKB_XI11.XI26.MM26_d
+ N_XI11.XI26.NET35_XI11.XI26.MM26_g N_VSS_XI11.XI26.MM26_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI24.MM26 N_XI11.XI24.CLKB_XI11.XI24.MM26_d
+ N_XI11.XI24.NET35_XI11.XI24.MM26_g N_VSS_XI11.XI24.MM26_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI27.MM26 N_XI11.XI27.CLKB_XI11.XI27.MM26_d
+ N_XI11.XI27.NET35_XI11.XI27.MM26_g N_VSS_XI11.XI27.MM26_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI22.MM26 N_XI11.XI22.CLKB_XI11.XI22.MM26_d
+ N_XI11.XI22.NET35_XI11.XI22.MM26_g N_VSS_XI11.XI22.MM26_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI21.MM26 N_XI11.XI21.CLKB_XI11.XI21.MM26_d
+ N_XI11.XI21.NET35_XI11.XI21.MM26_g N_VSS_XI11.XI21.MM26_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI23.MM26 N_XI11.XI23.CLKB_XI11.XI23.MM26_d
+ N_XI11.XI23.NET35_XI11.XI23.MM26_g N_VSS_XI11.XI23.MM26_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI19.MM26 N_XI11.XI19.CLKB_XI11.XI19.MM26_d
+ N_XI11.XI19.NET35_XI11.XI19.MM26_g N_VSS_XI11.XI19.MM26_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI20.MM26 N_XI11.XI20.CLKB_XI11.XI20.MM26_d
+ N_XI11.XI20.NET35_XI11.XI20.MM26_g N_VSS_XI11.XI20.MM26_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI18.MM26 N_XI11.XI18.CLKB_XI11.XI18.MM26_d
+ N_XI11.XI18.NET35_XI11.XI18.MM26_g N_VSS_XI11.XI18.MM26_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI17.MM26 N_XI11.XI17.CLKB_XI11.XI17.MM26_d
+ N_XI11.XI17.NET35_XI11.XI17.MM26_g N_VSS_XI11.XI17.MM26_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI0.MM26 N_XI11.XI0.CLKB_XI11.XI0.MM26_d N_XI11.XI0.NET35_XI11.XI0.MM26_g
+ N_VSS_XI11.XI0.MM26_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI11.XI30.MM19 N_XI11.XI30.NET27_XI11.XI30.MM19_d N_NET452_XI11.XI30.MM19_g
+ N_VSS_XI11.XI30.MM19_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI11.XI29.MM19 N_XI11.XI29.NET27_XI11.XI29.MM19_d N_NET453_XI11.XI29.MM19_g
+ N_VSS_XI11.XI29.MM19_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI11.XI31.MM19 N_XI11.XI31.NET27_XI11.XI31.MM19_d N_NET454_XI11.XI31.MM19_g
+ N_VSS_XI11.XI31.MM19_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI11.XI28.MM19 N_XI11.XI28.NET27_XI11.XI28.MM19_d N_NET455_XI11.XI28.MM19_g
+ N_VSS_XI11.XI28.MM19_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI11.XI25.MM19 N_XI11.XI25.NET27_XI11.XI25.MM19_d N_NET456_XI11.XI25.MM19_g
+ N_VSS_XI11.XI25.MM19_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI11.XI26.MM19 N_XI11.XI26.NET27_XI11.XI26.MM19_d N_NET457_XI11.XI26.MM19_g
+ N_VSS_XI11.XI26.MM19_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI11.XI24.MM19 N_XI11.XI24.NET27_XI11.XI24.MM19_d N_NET458_XI11.XI24.MM19_g
+ N_VSS_XI11.XI24.MM19_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI11.XI27.MM19 N_XI11.XI27.NET27_XI11.XI27.MM19_d N_NET459_XI11.XI27.MM19_g
+ N_VSS_XI11.XI27.MM19_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI11.XI22.MM19 N_XI11.XI22.NET27_XI11.XI22.MM19_d N_NET460_XI11.XI22.MM19_g
+ N_VSS_XI11.XI22.MM19_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI11.XI21.MM19 N_XI11.XI21.NET27_XI11.XI21.MM19_d N_NET461_XI11.XI21.MM19_g
+ N_VSS_XI11.XI21.MM19_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI11.XI23.MM19 N_XI11.XI23.NET27_XI11.XI23.MM19_d N_NET462_XI11.XI23.MM19_g
+ N_VSS_XI11.XI23.MM19_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI11.XI19.MM19 N_XI11.XI19.NET27_XI11.XI19.MM19_d N_NET463_XI11.XI19.MM19_g
+ N_VSS_XI11.XI19.MM19_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI11.XI20.MM19 N_XI11.XI20.NET27_XI11.XI20.MM19_d N_NET464_XI11.XI20.MM19_g
+ N_VSS_XI11.XI20.MM19_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI11.XI18.MM19 N_XI11.XI18.NET27_XI11.XI18.MM19_d N_NET465_XI11.XI18.MM19_g
+ N_VSS_XI11.XI18.MM19_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI11.XI17.MM19 N_XI11.XI17.NET27_XI11.XI17.MM19_d N_NET466_XI11.XI17.MM19_g
+ N_VSS_XI11.XI17.MM19_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI11.XI0.MM19 N_XI11.XI0.NET27_XI11.XI0.MM19_d N_NET467_XI11.XI0.MM19_g
+ N_VSS_XI11.XI0.MM19_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI11.XI30.MM18 N_XI11.XI30.NET31_XI11.XI30.MM18_d
+ N_XI11.XI30.NET27_XI11.XI30.MM18_g N_VSS_XI11.XI30.MM18_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI29.MM18 N_XI11.XI29.NET31_XI11.XI29.MM18_d
+ N_XI11.XI29.NET27_XI11.XI29.MM18_g N_VSS_XI11.XI29.MM18_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI31.MM18 N_XI11.XI31.NET31_XI11.XI31.MM18_d
+ N_XI11.XI31.NET27_XI11.XI31.MM18_g N_VSS_XI11.XI31.MM18_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI28.MM18 N_XI11.XI28.NET31_XI11.XI28.MM18_d
+ N_XI11.XI28.NET27_XI11.XI28.MM18_g N_VSS_XI11.XI28.MM18_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI25.MM18 N_XI11.XI25.NET31_XI11.XI25.MM18_d
+ N_XI11.XI25.NET27_XI11.XI25.MM18_g N_VSS_XI11.XI25.MM18_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI26.MM18 N_XI11.XI26.NET31_XI11.XI26.MM18_d
+ N_XI11.XI26.NET27_XI11.XI26.MM18_g N_VSS_XI11.XI26.MM18_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI24.MM18 N_XI11.XI24.NET31_XI11.XI24.MM18_d
+ N_XI11.XI24.NET27_XI11.XI24.MM18_g N_VSS_XI11.XI24.MM18_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI27.MM18 N_XI11.XI27.NET31_XI11.XI27.MM18_d
+ N_XI11.XI27.NET27_XI11.XI27.MM18_g N_VSS_XI11.XI27.MM18_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI22.MM18 N_XI11.XI22.NET31_XI11.XI22.MM18_d
+ N_XI11.XI22.NET27_XI11.XI22.MM18_g N_VSS_XI11.XI22.MM18_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI21.MM18 N_XI11.XI21.NET31_XI11.XI21.MM18_d
+ N_XI11.XI21.NET27_XI11.XI21.MM18_g N_VSS_XI11.XI21.MM18_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI23.MM18 N_XI11.XI23.NET31_XI11.XI23.MM18_d
+ N_XI11.XI23.NET27_XI11.XI23.MM18_g N_VSS_XI11.XI23.MM18_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI19.MM18 N_XI11.XI19.NET31_XI11.XI19.MM18_d
+ N_XI11.XI19.NET27_XI11.XI19.MM18_g N_VSS_XI11.XI19.MM18_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI20.MM18 N_XI11.XI20.NET31_XI11.XI20.MM18_d
+ N_XI11.XI20.NET27_XI11.XI20.MM18_g N_VSS_XI11.XI20.MM18_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI18.MM18 N_XI11.XI18.NET31_XI11.XI18.MM18_d
+ N_XI11.XI18.NET27_XI11.XI18.MM18_g N_VSS_XI11.XI18.MM18_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI17.MM18 N_XI11.XI17.NET31_XI11.XI17.MM18_d
+ N_XI11.XI17.NET27_XI11.XI17.MM18_g N_VSS_XI11.XI17.MM18_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI0.MM18 N_XI11.XI0.NET31_XI11.XI0.MM18_d N_XI11.XI0.NET27_XI11.XI0.MM18_g
+ N_VSS_XI11.XI0.MM18_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI11.XI30.MM28 N_XI11.XI30.NET31_XI11.XI30.MM28_d
+ N_XI11.XI30.CLKB_XI11.XI30.MM28_g N_XI11.XI30.NET58_XI11.XI30.MM28_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI29.MM28 N_XI11.XI29.NET31_XI11.XI29.MM28_d
+ N_XI11.XI29.CLKB_XI11.XI29.MM28_g N_XI11.XI29.NET58_XI11.XI29.MM28_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI31.MM28 N_XI11.XI31.NET31_XI11.XI31.MM28_d
+ N_XI11.XI31.CLKB_XI11.XI31.MM28_g N_XI11.XI31.NET58_XI11.XI31.MM28_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI28.MM28 N_XI11.XI28.NET31_XI11.XI28.MM28_d
+ N_XI11.XI28.CLKB_XI11.XI28.MM28_g N_XI11.XI28.NET58_XI11.XI28.MM28_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI25.MM28 N_XI11.XI25.NET31_XI11.XI25.MM28_d
+ N_XI11.XI25.CLKB_XI11.XI25.MM28_g N_XI11.XI25.NET58_XI11.XI25.MM28_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI26.MM28 N_XI11.XI26.NET31_XI11.XI26.MM28_d
+ N_XI11.XI26.CLKB_XI11.XI26.MM28_g N_XI11.XI26.NET58_XI11.XI26.MM28_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI24.MM28 N_XI11.XI24.NET31_XI11.XI24.MM28_d
+ N_XI11.XI24.CLKB_XI11.XI24.MM28_g N_XI11.XI24.NET58_XI11.XI24.MM28_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI27.MM28 N_XI11.XI27.NET31_XI11.XI27.MM28_d
+ N_XI11.XI27.CLKB_XI11.XI27.MM28_g N_XI11.XI27.NET58_XI11.XI27.MM28_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI22.MM28 N_XI11.XI22.NET31_XI11.XI22.MM28_d
+ N_XI11.XI22.CLKB_XI11.XI22.MM28_g N_XI11.XI22.NET58_XI11.XI22.MM28_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI21.MM28 N_XI11.XI21.NET31_XI11.XI21.MM28_d
+ N_XI11.XI21.CLKB_XI11.XI21.MM28_g N_XI11.XI21.NET58_XI11.XI21.MM28_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI23.MM28 N_XI11.XI23.NET31_XI11.XI23.MM28_d
+ N_XI11.XI23.CLKB_XI11.XI23.MM28_g N_XI11.XI23.NET58_XI11.XI23.MM28_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI19.MM28 N_XI11.XI19.NET31_XI11.XI19.MM28_d
+ N_XI11.XI19.CLKB_XI11.XI19.MM28_g N_XI11.XI19.NET58_XI11.XI19.MM28_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI20.MM28 N_XI11.XI20.NET31_XI11.XI20.MM28_d
+ N_XI11.XI20.CLKB_XI11.XI20.MM28_g N_XI11.XI20.NET58_XI11.XI20.MM28_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI18.MM28 N_XI11.XI18.NET31_XI11.XI18.MM28_d
+ N_XI11.XI18.CLKB_XI11.XI18.MM28_g N_XI11.XI18.NET58_XI11.XI18.MM28_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI17.MM28 N_XI11.XI17.NET31_XI11.XI17.MM28_d
+ N_XI11.XI17.CLKB_XI11.XI17.MM28_g N_XI11.XI17.NET58_XI11.XI17.MM28_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI0.MM28 N_XI11.XI0.NET31_XI11.XI0.MM28_d N_XI11.XI0.CLKB_XI11.XI0.MM28_g
+ N_XI11.XI0.NET58_XI11.XI0.MM28_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI11.XI30.MM6 N_XI11.XI30.NET15_XI11.XI30.MM6_d
+ N_XI11.XI30.NET58_XI11.XI30.MM6_g N_VSS_XI11.XI30.MM6_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI29.MM6 N_XI11.XI29.NET15_XI11.XI29.MM6_d
+ N_XI11.XI29.NET58_XI11.XI29.MM6_g N_VSS_XI11.XI29.MM6_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI31.MM6 N_XI11.XI31.NET15_XI11.XI31.MM6_d
+ N_XI11.XI31.NET58_XI11.XI31.MM6_g N_VSS_XI11.XI31.MM6_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI28.MM6 N_XI11.XI28.NET15_XI11.XI28.MM6_d
+ N_XI11.XI28.NET58_XI11.XI28.MM6_g N_VSS_XI11.XI28.MM6_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI25.MM6 N_XI11.XI25.NET15_XI11.XI25.MM6_d
+ N_XI11.XI25.NET58_XI11.XI25.MM6_g N_VSS_XI11.XI25.MM6_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI26.MM6 N_XI11.XI26.NET15_XI11.XI26.MM6_d
+ N_XI11.XI26.NET58_XI11.XI26.MM6_g N_VSS_XI11.XI26.MM6_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI24.MM6 N_XI11.XI24.NET15_XI11.XI24.MM6_d
+ N_XI11.XI24.NET58_XI11.XI24.MM6_g N_VSS_XI11.XI24.MM6_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI27.MM6 N_XI11.XI27.NET15_XI11.XI27.MM6_d
+ N_XI11.XI27.NET58_XI11.XI27.MM6_g N_VSS_XI11.XI27.MM6_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI22.MM6 N_XI11.XI22.NET15_XI11.XI22.MM6_d
+ N_XI11.XI22.NET58_XI11.XI22.MM6_g N_VSS_XI11.XI22.MM6_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI21.MM6 N_XI11.XI21.NET15_XI11.XI21.MM6_d
+ N_XI11.XI21.NET58_XI11.XI21.MM6_g N_VSS_XI11.XI21.MM6_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI23.MM6 N_XI11.XI23.NET15_XI11.XI23.MM6_d
+ N_XI11.XI23.NET58_XI11.XI23.MM6_g N_VSS_XI11.XI23.MM6_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI19.MM6 N_XI11.XI19.NET15_XI11.XI19.MM6_d
+ N_XI11.XI19.NET58_XI11.XI19.MM6_g N_VSS_XI11.XI19.MM6_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI20.MM6 N_XI11.XI20.NET15_XI11.XI20.MM6_d
+ N_XI11.XI20.NET58_XI11.XI20.MM6_g N_VSS_XI11.XI20.MM6_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI18.MM6 N_XI11.XI18.NET15_XI11.XI18.MM6_d
+ N_XI11.XI18.NET58_XI11.XI18.MM6_g N_VSS_XI11.XI18.MM6_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI17.MM6 N_XI11.XI17.NET15_XI11.XI17.MM6_d
+ N_XI11.XI17.NET58_XI11.XI17.MM6_g N_VSS_XI11.XI17.MM6_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI0.MM6 N_XI11.XI0.NET15_XI11.XI0.MM6_d N_XI11.XI0.NET58_XI11.XI0.MM6_g
+ N_VSS_XI11.XI0.MM6_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI11.XI30.MM0 N_XI11.XI30.NET54_XI11.XI30.MM0_d
+ N_XI11.XI30.NET15_XI11.XI30.MM0_g N_VSS_XI11.XI30.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI29.MM0 N_XI11.XI29.NET54_XI11.XI29.MM0_d
+ N_XI11.XI29.NET15_XI11.XI29.MM0_g N_VSS_XI11.XI29.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI31.MM0 N_XI11.XI31.NET54_XI11.XI31.MM0_d
+ N_XI11.XI31.NET15_XI11.XI31.MM0_g N_VSS_XI11.XI31.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI28.MM0 N_XI11.XI28.NET54_XI11.XI28.MM0_d
+ N_XI11.XI28.NET15_XI11.XI28.MM0_g N_VSS_XI11.XI28.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI25.MM0 N_XI11.XI25.NET54_XI11.XI25.MM0_d
+ N_XI11.XI25.NET15_XI11.XI25.MM0_g N_VSS_XI11.XI25.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI26.MM0 N_XI11.XI26.NET54_XI11.XI26.MM0_d
+ N_XI11.XI26.NET15_XI11.XI26.MM0_g N_VSS_XI11.XI26.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI24.MM0 N_XI11.XI24.NET54_XI11.XI24.MM0_d
+ N_XI11.XI24.NET15_XI11.XI24.MM0_g N_VSS_XI11.XI24.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI27.MM0 N_XI11.XI27.NET54_XI11.XI27.MM0_d
+ N_XI11.XI27.NET15_XI11.XI27.MM0_g N_VSS_XI11.XI27.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI22.MM0 N_XI11.XI22.NET54_XI11.XI22.MM0_d
+ N_XI11.XI22.NET15_XI11.XI22.MM0_g N_VSS_XI11.XI22.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI21.MM0 N_XI11.XI21.NET54_XI11.XI21.MM0_d
+ N_XI11.XI21.NET15_XI11.XI21.MM0_g N_VSS_XI11.XI21.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI23.MM0 N_XI11.XI23.NET54_XI11.XI23.MM0_d
+ N_XI11.XI23.NET15_XI11.XI23.MM0_g N_VSS_XI11.XI23.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI19.MM0 N_XI11.XI19.NET54_XI11.XI19.MM0_d
+ N_XI11.XI19.NET15_XI11.XI19.MM0_g N_VSS_XI11.XI19.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI20.MM0 N_XI11.XI20.NET54_XI11.XI20.MM0_d
+ N_XI11.XI20.NET15_XI11.XI20.MM0_g N_VSS_XI11.XI20.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI18.MM0 N_XI11.XI18.NET54_XI11.XI18.MM0_d
+ N_XI11.XI18.NET15_XI11.XI18.MM0_g N_VSS_XI11.XI18.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI17.MM0 N_XI11.XI17.NET54_XI11.XI17.MM0_d
+ N_XI11.XI17.NET15_XI11.XI17.MM0_g N_VSS_XI11.XI17.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI0.MM0 N_XI11.XI0.NET54_XI11.XI0.MM0_d N_XI11.XI0.NET15_XI11.XI0.MM0_g
+ N_VSS_XI11.XI0.MM0_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI11.XI30.MM36 N_XI11.XI30.NET58_XI11.XI30.MM36_d
+ N_XI11.XI30.NET35_XI11.XI30.MM36_g N_XI11.XI30.NET54_XI11.XI30.MM36_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI29.MM36 N_XI11.XI29.NET58_XI11.XI29.MM36_d
+ N_XI11.XI29.NET35_XI11.XI29.MM36_g N_XI11.XI29.NET54_XI11.XI29.MM36_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI31.MM36 N_XI11.XI31.NET58_XI11.XI31.MM36_d
+ N_XI11.XI31.NET35_XI11.XI31.MM36_g N_XI11.XI31.NET54_XI11.XI31.MM36_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI28.MM36 N_XI11.XI28.NET58_XI11.XI28.MM36_d
+ N_XI11.XI28.NET35_XI11.XI28.MM36_g N_XI11.XI28.NET54_XI11.XI28.MM36_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI25.MM36 N_XI11.XI25.NET58_XI11.XI25.MM36_d
+ N_XI11.XI25.NET35_XI11.XI25.MM36_g N_XI11.XI25.NET54_XI11.XI25.MM36_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI26.MM36 N_XI11.XI26.NET58_XI11.XI26.MM36_d
+ N_XI11.XI26.NET35_XI11.XI26.MM36_g N_XI11.XI26.NET54_XI11.XI26.MM36_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI24.MM36 N_XI11.XI24.NET58_XI11.XI24.MM36_d
+ N_XI11.XI24.NET35_XI11.XI24.MM36_g N_XI11.XI24.NET54_XI11.XI24.MM36_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI27.MM36 N_XI11.XI27.NET58_XI11.XI27.MM36_d
+ N_XI11.XI27.NET35_XI11.XI27.MM36_g N_XI11.XI27.NET54_XI11.XI27.MM36_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI22.MM36 N_XI11.XI22.NET58_XI11.XI22.MM36_d
+ N_XI11.XI22.NET35_XI11.XI22.MM36_g N_XI11.XI22.NET54_XI11.XI22.MM36_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI21.MM36 N_XI11.XI21.NET58_XI11.XI21.MM36_d
+ N_XI11.XI21.NET35_XI11.XI21.MM36_g N_XI11.XI21.NET54_XI11.XI21.MM36_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI23.MM36 N_XI11.XI23.NET58_XI11.XI23.MM36_d
+ N_XI11.XI23.NET35_XI11.XI23.MM36_g N_XI11.XI23.NET54_XI11.XI23.MM36_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI19.MM36 N_XI11.XI19.NET58_XI11.XI19.MM36_d
+ N_XI11.XI19.NET35_XI11.XI19.MM36_g N_XI11.XI19.NET54_XI11.XI19.MM36_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI20.MM36 N_XI11.XI20.NET58_XI11.XI20.MM36_d
+ N_XI11.XI20.NET35_XI11.XI20.MM36_g N_XI11.XI20.NET54_XI11.XI20.MM36_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI18.MM36 N_XI11.XI18.NET58_XI11.XI18.MM36_d
+ N_XI11.XI18.NET35_XI11.XI18.MM36_g N_XI11.XI18.NET54_XI11.XI18.MM36_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI17.MM36 N_XI11.XI17.NET58_XI11.XI17.MM36_d
+ N_XI11.XI17.NET35_XI11.XI17.MM36_g N_XI11.XI17.NET54_XI11.XI17.MM36_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI0.MM36 N_XI11.XI0.NET58_XI11.XI0.MM36_d N_XI11.XI0.NET35_XI11.XI0.MM36_g
+ N_XI11.XI0.NET54_XI11.XI0.MM36_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI11.XI30.MM38 N_XI11.XI30.NET15_XI11.XI30.MM38_d
+ N_XI11.XI30.NET35_XI11.XI30.MM38_g N_XI11.XI30.NET14_XI11.XI30.MM38_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI29.MM38 N_XI11.XI29.NET15_XI11.XI29.MM38_d
+ N_XI11.XI29.NET35_XI11.XI29.MM38_g N_XI11.XI29.NET14_XI11.XI29.MM38_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI31.MM38 N_XI11.XI31.NET15_XI11.XI31.MM38_d
+ N_XI11.XI31.NET35_XI11.XI31.MM38_g N_XI11.XI31.NET14_XI11.XI31.MM38_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI28.MM38 N_XI11.XI28.NET15_XI11.XI28.MM38_d
+ N_XI11.XI28.NET35_XI11.XI28.MM38_g N_XI11.XI28.NET14_XI11.XI28.MM38_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI25.MM38 N_XI11.XI25.NET15_XI11.XI25.MM38_d
+ N_XI11.XI25.NET35_XI11.XI25.MM38_g N_XI11.XI25.NET14_XI11.XI25.MM38_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI26.MM38 N_XI11.XI26.NET15_XI11.XI26.MM38_d
+ N_XI11.XI26.NET35_XI11.XI26.MM38_g N_XI11.XI26.NET14_XI11.XI26.MM38_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI24.MM38 N_XI11.XI24.NET15_XI11.XI24.MM38_d
+ N_XI11.XI24.NET35_XI11.XI24.MM38_g N_XI11.XI24.NET14_XI11.XI24.MM38_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI27.MM38 N_XI11.XI27.NET15_XI11.XI27.MM38_d
+ N_XI11.XI27.NET35_XI11.XI27.MM38_g N_XI11.XI27.NET14_XI11.XI27.MM38_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI22.MM38 N_XI11.XI22.NET15_XI11.XI22.MM38_d
+ N_XI11.XI22.NET35_XI11.XI22.MM38_g N_XI11.XI22.NET14_XI11.XI22.MM38_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI21.MM38 N_XI11.XI21.NET15_XI11.XI21.MM38_d
+ N_XI11.XI21.NET35_XI11.XI21.MM38_g N_XI11.XI21.NET14_XI11.XI21.MM38_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI23.MM38 N_XI11.XI23.NET15_XI11.XI23.MM38_d
+ N_XI11.XI23.NET35_XI11.XI23.MM38_g N_XI11.XI23.NET14_XI11.XI23.MM38_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI19.MM38 N_XI11.XI19.NET15_XI11.XI19.MM38_d
+ N_XI11.XI19.NET35_XI11.XI19.MM38_g N_XI11.XI19.NET14_XI11.XI19.MM38_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI20.MM38 N_XI11.XI20.NET15_XI11.XI20.MM38_d
+ N_XI11.XI20.NET35_XI11.XI20.MM38_g N_XI11.XI20.NET14_XI11.XI20.MM38_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI18.MM38 N_XI11.XI18.NET15_XI11.XI18.MM38_d
+ N_XI11.XI18.NET35_XI11.XI18.MM38_g N_XI11.XI18.NET14_XI11.XI18.MM38_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI17.MM38 N_XI11.XI17.NET15_XI11.XI17.MM38_d
+ N_XI11.XI17.NET35_XI11.XI17.MM38_g N_XI11.XI17.NET14_XI11.XI17.MM38_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI0.MM38 N_XI11.XI0.NET15_XI11.XI0.MM38_d N_XI11.XI0.NET35_XI11.XI0.MM38_g
+ N_XI11.XI0.NET14_XI11.XI0.MM38_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI11.XI30.MM15 N_ACC15_XI11.XI30.MM15_d N_XI11.XI30.NET14_XI11.XI30.MM15_g
+ N_VSS_XI11.XI30.MM15_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI11.XI29.MM15 N_ACC14_XI11.XI29.MM15_d N_XI11.XI29.NET14_XI11.XI29.MM15_g
+ N_VSS_XI11.XI29.MM15_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI11.XI31.MM15 N_ACC13_XI11.XI31.MM15_d N_XI11.XI31.NET14_XI11.XI31.MM15_g
+ N_VSS_XI11.XI31.MM15_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI11.XI28.MM15 N_ACC12_XI11.XI28.MM15_d N_XI11.XI28.NET14_XI11.XI28.MM15_g
+ N_VSS_XI11.XI28.MM15_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI11.XI25.MM15 N_ACC11_XI11.XI25.MM15_d N_XI11.XI25.NET14_XI11.XI25.MM15_g
+ N_VSS_XI11.XI25.MM15_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI11.XI26.MM15 N_ACC10_XI11.XI26.MM15_d N_XI11.XI26.NET14_XI11.XI26.MM15_g
+ N_VSS_XI11.XI26.MM15_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI11.XI24.MM15 N_ACC9_XI11.XI24.MM15_d N_XI11.XI24.NET14_XI11.XI24.MM15_g
+ N_VSS_XI11.XI24.MM15_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI11.XI27.MM15 N_ACC8_XI11.XI27.MM15_d N_XI11.XI27.NET14_XI11.XI27.MM15_g
+ N_VSS_XI11.XI27.MM15_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI11.XI22.MM15 N_ACC7_XI11.XI22.MM15_d N_XI11.XI22.NET14_XI11.XI22.MM15_g
+ N_VSS_XI11.XI22.MM15_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI11.XI21.MM15 N_ACC6_XI11.XI21.MM15_d N_XI11.XI21.NET14_XI11.XI21.MM15_g
+ N_VSS_XI11.XI21.MM15_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI11.XI23.MM15 N_ACC5_XI11.XI23.MM15_d N_XI11.XI23.NET14_XI11.XI23.MM15_g
+ N_VSS_XI11.XI23.MM15_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI11.XI19.MM15 N_ACC4_XI11.XI19.MM15_d N_XI11.XI19.NET14_XI11.XI19.MM15_g
+ N_VSS_XI11.XI19.MM15_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI11.XI20.MM15 N_ACC3_XI11.XI20.MM15_d N_XI11.XI20.NET14_XI11.XI20.MM15_g
+ N_VSS_XI11.XI20.MM15_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI11.XI18.MM15 N_ACC2_XI11.XI18.MM15_d N_XI11.XI18.NET14_XI11.XI18.MM15_g
+ N_VSS_XI11.XI18.MM15_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI11.XI17.MM15 N_ACC1_XI11.XI17.MM15_d N_XI11.XI17.NET14_XI11.XI17.MM15_g
+ N_VSS_XI11.XI17.MM15_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI11.XI0.MM15 N_ACC0_XI11.XI0.MM15_d N_XI11.XI0.NET14_XI11.XI0.MM15_g
+ N_VSS_XI11.XI0.MM15_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI11.XI30.MM16 N_XI11.BAR_Q16_XI11.XI30.MM16_d N_ACC15_XI11.XI30.MM16_g
+ N_VSS_XI11.XI30.MM16_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI11.XI29.MM16 N_XI11.BAR_Q15_XI11.XI29.MM16_d N_ACC14_XI11.XI29.MM16_g
+ N_VSS_XI11.XI29.MM16_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI11.XI31.MM16 N_XI11.BAR_Q14_XI11.XI31.MM16_d N_ACC13_XI11.XI31.MM16_g
+ N_VSS_XI11.XI31.MM16_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI11.XI28.MM16 N_XI11.BAR_Q13_XI11.XI28.MM16_d N_ACC12_XI11.XI28.MM16_g
+ N_VSS_XI11.XI28.MM16_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI11.XI25.MM16 N_XI11.BAR_Q12_XI11.XI25.MM16_d N_ACC11_XI11.XI25.MM16_g
+ N_VSS_XI11.XI25.MM16_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI11.XI26.MM16 N_XI11.BAR_Q11_XI11.XI26.MM16_d N_ACC10_XI11.XI26.MM16_g
+ N_VSS_XI11.XI26.MM16_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI11.XI24.MM16 N_XI11.BAR_Q10_XI11.XI24.MM16_d N_ACC9_XI11.XI24.MM16_g
+ N_VSS_XI11.XI24.MM16_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI11.XI27.MM16 N_XI11.BAR_Q9_XI11.XI27.MM16_d N_ACC8_XI11.XI27.MM16_g
+ N_VSS_XI11.XI27.MM16_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI11.XI22.MM16 N_XI11.BAR_Q8_XI11.XI22.MM16_d N_ACC7_XI11.XI22.MM16_g
+ N_VSS_XI11.XI22.MM16_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI11.XI21.MM16 N_XI11.BAR_Q7_XI11.XI21.MM16_d N_ACC6_XI11.XI21.MM16_g
+ N_VSS_XI11.XI21.MM16_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI11.XI23.MM16 N_XI11.BAR_Q6_XI11.XI23.MM16_d N_ACC5_XI11.XI23.MM16_g
+ N_VSS_XI11.XI23.MM16_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI11.XI19.MM16 N_XI11.BAR_Q5_XI11.XI19.MM16_d N_ACC4_XI11.XI19.MM16_g
+ N_VSS_XI11.XI19.MM16_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI11.XI20.MM16 N_XI11.BAR_Q4_XI11.XI20.MM16_d N_ACC3_XI11.XI20.MM16_g
+ N_VSS_XI11.XI20.MM16_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI11.XI18.MM16 N_XI11.BAR_Q3_XI11.XI18.MM16_d N_ACC2_XI11.XI18.MM16_g
+ N_VSS_XI11.XI18.MM16_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI11.XI17.MM16 N_XI11.BAR_Q2_XI11.XI17.MM16_d N_ACC1_XI11.XI17.MM16_g
+ N_VSS_XI11.XI17.MM16_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI11.XI0.MM16 N_XI11.BAR_Q1_XI11.XI0.MM16_d N_ACC0_XI11.XI0.MM16_g
+ N_VSS_XI11.XI0.MM16_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI11.XI30.MM40 N_XI11.XI30.NET14_XI11.XI30.MM40_d
+ N_XI11.XI30.CLKB_XI11.XI30.MM40_g N_XI11.BAR_Q16_XI11.XI30.MM40_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI29.MM40 N_XI11.XI29.NET14_XI11.XI29.MM40_d
+ N_XI11.XI29.CLKB_XI11.XI29.MM40_g N_XI11.BAR_Q15_XI11.XI29.MM40_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI31.MM40 N_XI11.XI31.NET14_XI11.XI31.MM40_d
+ N_XI11.XI31.CLKB_XI11.XI31.MM40_g N_XI11.BAR_Q14_XI11.XI31.MM40_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI28.MM40 N_XI11.XI28.NET14_XI11.XI28.MM40_d
+ N_XI11.XI28.CLKB_XI11.XI28.MM40_g N_XI11.BAR_Q13_XI11.XI28.MM40_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI25.MM40 N_XI11.XI25.NET14_XI11.XI25.MM40_d
+ N_XI11.XI25.CLKB_XI11.XI25.MM40_g N_XI11.BAR_Q12_XI11.XI25.MM40_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI26.MM40 N_XI11.XI26.NET14_XI11.XI26.MM40_d
+ N_XI11.XI26.CLKB_XI11.XI26.MM40_g N_XI11.BAR_Q11_XI11.XI26.MM40_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI24.MM40 N_XI11.XI24.NET14_XI11.XI24.MM40_d
+ N_XI11.XI24.CLKB_XI11.XI24.MM40_g N_XI11.BAR_Q10_XI11.XI24.MM40_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI27.MM40 N_XI11.XI27.NET14_XI11.XI27.MM40_d
+ N_XI11.XI27.CLKB_XI11.XI27.MM40_g N_XI11.BAR_Q9_XI11.XI27.MM40_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI22.MM40 N_XI11.XI22.NET14_XI11.XI22.MM40_d
+ N_XI11.XI22.CLKB_XI11.XI22.MM40_g N_XI11.BAR_Q8_XI11.XI22.MM40_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI21.MM40 N_XI11.XI21.NET14_XI11.XI21.MM40_d
+ N_XI11.XI21.CLKB_XI11.XI21.MM40_g N_XI11.BAR_Q7_XI11.XI21.MM40_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI23.MM40 N_XI11.XI23.NET14_XI11.XI23.MM40_d
+ N_XI11.XI23.CLKB_XI11.XI23.MM40_g N_XI11.BAR_Q6_XI11.XI23.MM40_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI19.MM40 N_XI11.XI19.NET14_XI11.XI19.MM40_d
+ N_XI11.XI19.CLKB_XI11.XI19.MM40_g N_XI11.BAR_Q5_XI11.XI19.MM40_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI20.MM40 N_XI11.XI20.NET14_XI11.XI20.MM40_d
+ N_XI11.XI20.CLKB_XI11.XI20.MM40_g N_XI11.BAR_Q4_XI11.XI20.MM40_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI18.MM40 N_XI11.XI18.NET14_XI11.XI18.MM40_d
+ N_XI11.XI18.CLKB_XI11.XI18.MM40_g N_XI11.BAR_Q3_XI11.XI18.MM40_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI17.MM40 N_XI11.XI17.NET14_XI11.XI17.MM40_d
+ N_XI11.XI17.CLKB_XI11.XI17.MM40_g N_XI11.BAR_Q2_XI11.XI17.MM40_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI11.XI0.MM40 N_XI11.XI0.NET14_XI11.XI0.MM40_d N_XI11.XI0.CLKB_XI11.XI0.MM40_g
+ N_XI11.BAR_Q1_XI11.XI0.MM40_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI20.XI11.MM2 N_NET594_XI20.XI11.MM2_d N_NET241_XI20.XI11.MM2_g
+ N_VSS_XI20.XI11.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI21.XI11.MM2 N_NET628_XI21.XI11.MM2_d N_NET241_XI21.XI11.MM2_g
+ N_VSS_XI21.XI11.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI20.XI12.MM2 N_NET595_XI20.XI12.MM2_d N_NET242_XI20.XI12.MM2_g
+ N_VSS_XI20.XI12.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI21.XI12.MM2 N_NET629_XI21.XI12.MM2_d N_NET242_XI21.XI12.MM2_g
+ N_VSS_XI21.XI12.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI20.XI10.MM2 N_NET596_XI20.XI10.MM2_d N_NET243_XI20.XI10.MM2_g
+ N_VSS_XI20.XI10.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI21.XI10.MM2 N_NET630_XI21.XI10.MM2_d N_NET243_XI21.XI10.MM2_g
+ N_VSS_XI21.XI10.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI20.XI9.MM2 N_NET597_XI20.XI9.MM2_d N_NET244_XI20.XI9.MM2_g
+ N_VSS_XI20.XI9.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI21.XI9.MM2 N_NET631_XI21.XI9.MM2_d N_NET244_XI21.XI9.MM2_g
+ N_VSS_XI21.XI9.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI20.XI14.MM2 N_NET598_XI20.XI14.MM2_d N_NET245_XI20.XI14.MM2_g
+ N_VSS_XI20.XI14.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI21.XI14.MM2 N_NET632_XI21.XI14.MM2_d N_NET245_XI21.XI14.MM2_g
+ N_VSS_XI21.XI14.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI20.XI13.MM2 N_NET599_XI20.XI13.MM2_d N_NET246_XI20.XI13.MM2_g
+ N_VSS_XI20.XI13.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI21.XI13.MM2 N_NET633_XI21.XI13.MM2_d N_NET246_XI21.XI13.MM2_g
+ N_VSS_XI21.XI13.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI20.XI15.MM2 N_NET600_XI20.XI15.MM2_d N_NET247_XI20.XI15.MM2_g
+ N_VSS_XI20.XI15.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI21.XI15.MM2 N_NET634_XI21.XI15.MM2_d N_NET247_XI21.XI15.MM2_g
+ N_VSS_XI21.XI15.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI20.XI6.MM2 N_NET601_XI20.XI6.MM2_d N_NET248_XI20.XI6.MM2_g
+ N_VSS_XI20.XI6.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI21.XI6.MM2 N_NET635_XI21.XI6.MM2_d N_NET248_XI21.XI6.MM2_g
+ N_VSS_XI21.XI6.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI20.XI5.MM2 N_NET602_XI20.XI5.MM2_d N_NET249_XI20.XI5.MM2_g
+ N_VSS_XI20.XI5.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI21.XI5.MM2 N_NET636_XI21.XI5.MM2_d N_NET249_XI21.XI5.MM2_g
+ N_VSS_XI21.XI5.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI20.XI7.MM2 N_NET603_XI20.XI7.MM2_d N_NET250_XI20.XI7.MM2_g
+ N_VSS_XI20.XI7.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI21.XI7.MM2 N_NET637_XI21.XI7.MM2_d N_NET250_XI21.XI7.MM2_g
+ N_VSS_XI21.XI7.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI20.XI8.MM2 N_NET604_XI20.XI8.MM2_d N_NET251_XI20.XI8.MM2_g
+ N_VSS_XI20.XI8.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI21.XI8.MM2 N_NET638_XI21.XI8.MM2_d N_NET251_XI21.XI8.MM2_g
+ N_VSS_XI21.XI8.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI20.XI3.MM2 N_NET605_XI20.XI3.MM2_d N_NET252_XI20.XI3.MM2_g
+ N_VSS_XI20.XI3.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI21.XI3.MM2 N_NET639_XI21.XI3.MM2_d N_NET252_XI21.XI3.MM2_g
+ N_VSS_XI21.XI3.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI20.XI4.MM2 N_NET606_XI20.XI4.MM2_d N_NET253_XI20.XI4.MM2_g
+ N_VSS_XI20.XI4.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI21.XI4.MM2 N_NET640_XI21.XI4.MM2_d N_NET253_XI21.XI4.MM2_g
+ N_VSS_XI21.XI4.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI20.XI2.MM2 N_NET607_XI20.XI2.MM2_d N_NET254_XI20.XI2.MM2_g
+ N_VSS_XI20.XI2.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI21.XI2.MM2 N_NET641_XI21.XI2.MM2_d N_NET254_XI21.XI2.MM2_g
+ N_VSS_XI21.XI2.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI20.XI1.MM2 N_NET608_XI20.XI1.MM2_d N_NET255_XI20.XI1.MM2_g
+ N_VSS_XI20.XI1.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI21.XI1.MM2 N_NET642_XI21.XI1.MM2_d N_NET255_XI21.XI1.MM2_g
+ N_VSS_XI21.XI1.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI20.XI0.MM2 N_NET609_XI20.XI0.MM2_d N_NET256_XI20.XI0.MM2_g
+ N_VSS_XI20.XI0.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI21.XI0.MM2 N_NET643_XI21.XI0.MM2_d N_NET256_XI21.XI0.MM2_g
+ N_VSS_XI21.XI0.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI0.XI134.XI9.MM2 N_XI0.XI134.NET43_XI0.XI134.XI9.MM2_d
+ N_NET594_XI0.XI134.XI9.MM2_g N_VSS_XI0.XI134.XI9.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI0.XI153.XI1.MM2 N_XI0.XI153.XI1.NET036_XI0.XI153.XI1.MM2_d
+ N_NET595_XI0.XI153.XI1.MM2_g N_VSS_XI0.XI153.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.85e-13 AS=2.45e-13
+ PD=7.4e-07 PS=1.48e-06
mXI0.XI154.XI1.MM2 N_XI0.XI154.XI1.NET036_XI0.XI154.XI1.MM2_d
+ N_NET596_XI0.XI154.XI1.MM2_g N_VSS_XI0.XI154.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.85e-13 AS=2.45e-13
+ PD=7.4e-07 PS=1.48e-06
mXI0.XI157.XI1.MM2 N_XI0.XI157.XI1.NET036_XI0.XI157.XI1.MM2_d
+ N_NET597_XI0.XI157.XI1.MM2_g N_VSS_XI0.XI157.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.85e-13 AS=2.45e-13
+ PD=7.4e-07 PS=1.48e-06
mXI0.XI156.XI1.MM2 N_XI0.XI156.XI1.NET036_XI0.XI156.XI1.MM2_d
+ N_NET598_XI0.XI156.XI1.MM2_g N_VSS_XI0.XI156.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.85e-13 AS=2.45e-13
+ PD=7.4e-07 PS=1.48e-06
mXI0.XI155.XI1.MM2 N_XI0.XI155.XI1.NET036_XI0.XI155.XI1.MM2_d
+ N_NET599_XI0.XI155.XI1.MM2_g N_VSS_XI0.XI155.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.85e-13 AS=2.45e-13
+ PD=7.4e-07 PS=1.48e-06
mXI0.XI133.XI1.MM2 N_XI0.XI133.XI1.NET036_XI0.XI133.XI1.MM2_d
+ N_NET600_XI0.XI133.XI1.MM2_g N_VSS_XI0.XI133.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.85e-13 AS=2.45e-13
+ PD=7.4e-07 PS=1.48e-06
mXI0.XI132.XI1.MM2 N_XI0.XI132.XI1.NET036_XI0.XI132.XI1.MM2_d
+ N_NET601_XI0.XI132.XI1.MM2_g N_VSS_XI0.XI132.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.85e-13 AS=2.45e-13
+ PD=7.4e-07 PS=1.48e-06
mXI0.XI131.XI1.MM2 N_XI0.XI131.XI1.NET036_XI0.XI131.XI1.MM2_d
+ N_NET602_XI0.XI131.XI1.MM2_g N_VSS_XI0.XI131.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.85e-13 AS=2.45e-13
+ PD=7.4e-07 PS=1.48e-06
mXI0.XI111.XI1.MM2 N_XI0.XI111.XI1.NET036_XI0.XI111.XI1.MM2_d
+ N_NET603_XI0.XI111.XI1.MM2_g N_VSS_XI0.XI111.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.85e-13 AS=2.45e-13
+ PD=7.4e-07 PS=1.48e-06
mXI0.XI110.XI1.MM2 N_XI0.XI110.XI1.NET036_XI0.XI110.XI1.MM2_d
+ N_NET604_XI0.XI110.XI1.MM2_g N_VSS_XI0.XI110.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.85e-13 AS=2.45e-13
+ PD=7.4e-07 PS=1.48e-06
mXI0.XI103.XI1.MM2 N_XI0.XI103.XI1.NET036_XI0.XI103.XI1.MM2_d
+ N_NET605_XI0.XI103.XI1.MM2_g N_VSS_XI0.XI103.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.85e-13 AS=2.45e-13
+ PD=7.4e-07 PS=1.48e-06
mXI0.XI102.XI1.MM2 N_XI0.XI102.XI1.NET036_XI0.XI102.XI1.MM2_d
+ N_NET606_XI0.XI102.XI1.MM2_g N_VSS_XI0.XI102.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.85e-13 AS=2.45e-13
+ PD=7.4e-07 PS=1.48e-06
mXI0.XI88.XI1.MM2 N_XI0.XI88.XI1.NET036_XI0.XI88.XI1.MM2_d
+ N_NET607_XI0.XI88.XI1.MM2_g N_VSS_XI0.XI88.XI1.MM2_s N_VSS_XI10.XI0.XI0.MM2_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.85e-13 AS=2.45e-13 PD=7.4e-07 PS=1.48e-06
mXI0.XI82.XI1.MM2 N_XI0.XI82.XI1.NET036_XI0.XI82.XI1.MM2_d
+ N_NET608_XI0.XI82.XI1.MM2_g N_VSS_XI0.XI82.XI1.MM2_s N_VSS_XI10.XI0.XI0.MM2_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.85e-13 AS=2.45e-13 PD=7.4e-07 PS=1.48e-06
mXI0.XI10.XI1.MM2 N_XI0.XI10.XI1.NET036_XI0.XI10.XI1.MM2_d
+ N_NET609_XI0.XI10.XI1.MM2_g N_VSS_XI0.XI10.XI1.MM2_s N_VSS_XI10.XI0.XI0.MM2_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.85e-13 AS=2.45e-13 PD=7.4e-07 PS=1.48e-06
mXI0.XI153.XI1.MM0 N_XI0.XI153.NET6_XI0.XI153.XI1.MM0_d
+ N_MIN14_XI0.XI153.XI1.MM0_g N_XI0.XI153.XI1.NET036_XI0.XI153.XI1.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=1.85e-13
+ PD=1.52e-06 PS=7.4e-07
mXI0.XI154.XI1.MM0 N_XI0.XI154.NET6_XI0.XI154.XI1.MM0_d
+ N_MIN13_XI0.XI154.XI1.MM0_g N_XI0.XI154.XI1.NET036_XI0.XI154.XI1.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=1.85e-13
+ PD=1.52e-06 PS=7.4e-07
mXI0.XI157.XI1.MM0 N_XI0.XI157.NET6_XI0.XI157.XI1.MM0_d
+ N_MIN12_XI0.XI157.XI1.MM0_g N_XI0.XI157.XI1.NET036_XI0.XI157.XI1.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=1.85e-13
+ PD=1.52e-06 PS=7.4e-07
mXI0.XI156.XI1.MM0 N_XI0.XI156.NET6_XI0.XI156.XI1.MM0_d
+ N_MIN11_XI0.XI156.XI1.MM0_g N_XI0.XI156.XI1.NET036_XI0.XI156.XI1.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=1.85e-13
+ PD=1.52e-06 PS=7.4e-07
mXI0.XI155.XI1.MM0 N_XI0.XI155.NET6_XI0.XI155.XI1.MM0_d
+ N_MIN10_XI0.XI155.XI1.MM0_g N_XI0.XI155.XI1.NET036_XI0.XI155.XI1.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=1.85e-13
+ PD=1.52e-06 PS=7.4e-07
mXI0.XI133.XI1.MM0 N_XI0.XI133.NET6_XI0.XI133.XI1.MM0_d
+ N_MIN9_XI0.XI133.XI1.MM0_g N_XI0.XI133.XI1.NET036_XI0.XI133.XI1.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=1.85e-13
+ PD=1.52e-06 PS=7.4e-07
mXI0.XI132.XI1.MM0 N_XI0.XI132.NET6_XI0.XI132.XI1.MM0_d
+ N_MIN8_XI0.XI132.XI1.MM0_g N_XI0.XI132.XI1.NET036_XI0.XI132.XI1.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=1.85e-13
+ PD=1.52e-06 PS=7.4e-07
mXI0.XI131.XI1.MM0 N_XI0.XI131.NET6_XI0.XI131.XI1.MM0_d
+ N_MIN7_XI0.XI131.XI1.MM0_g N_XI0.XI131.XI1.NET036_XI0.XI131.XI1.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=1.85e-13
+ PD=1.52e-06 PS=7.4e-07
mXI0.XI111.XI1.MM0 N_XI0.XI111.NET6_XI0.XI111.XI1.MM0_d
+ N_MIN6_XI0.XI111.XI1.MM0_g N_XI0.XI111.XI1.NET036_XI0.XI111.XI1.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=1.85e-13
+ PD=1.52e-06 PS=7.4e-07
mXI0.XI110.XI1.MM0 N_XI0.XI110.NET6_XI0.XI110.XI1.MM0_d
+ N_MIN5_XI0.XI110.XI1.MM0_g N_XI0.XI110.XI1.NET036_XI0.XI110.XI1.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=1.85e-13
+ PD=1.52e-06 PS=7.4e-07
mXI0.XI103.XI1.MM0 N_XI0.XI103.NET6_XI0.XI103.XI1.MM0_d
+ N_MIN4_XI0.XI103.XI1.MM0_g N_XI0.XI103.XI1.NET036_XI0.XI103.XI1.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=1.85e-13
+ PD=1.52e-06 PS=7.4e-07
mXI0.XI102.XI1.MM0 N_XI0.XI102.NET6_XI0.XI102.XI1.MM0_d
+ N_MIN3_XI0.XI102.XI1.MM0_g N_XI0.XI102.XI1.NET036_XI0.XI102.XI1.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=1.85e-13
+ PD=1.52e-06 PS=7.4e-07
mXI0.XI88.XI1.MM0 N_XI0.XI88.NET6_XI0.XI88.XI1.MM0_d N_MIN2_XI0.XI88.XI1.MM0_g
+ N_XI0.XI88.XI1.NET036_XI0.XI88.XI1.MM0_s N_VSS_XI10.XI0.XI0.MM2_b N_18
+ L=1.8e-07 W=5e-07 AD=2.55e-13 AS=1.85e-13 PD=1.52e-06 PS=7.4e-07
mXI0.XI82.XI1.MM0 N_XI0.XI82.NET6_XI0.XI82.XI1.MM0_d N_MIN1_XI0.XI82.XI1.MM0_g
+ N_XI0.XI82.XI1.NET036_XI0.XI82.XI1.MM0_s N_VSS_XI10.XI0.XI0.MM2_b N_18
+ L=1.8e-07 W=5e-07 AD=2.55e-13 AS=1.85e-13 PD=1.52e-06 PS=7.4e-07
mXI0.XI10.XI1.MM0 N_XI0.XI10.NET6_XI0.XI10.XI1.MM0_d N_MIN0_XI0.XI10.XI1.MM0_g
+ N_XI0.XI10.XI1.NET036_XI0.XI10.XI1.MM0_s N_VSS_XI10.XI0.XI0.MM2_b N_18
+ L=1.8e-07 W=5e-07 AD=2.55e-13 AS=1.85e-13 PD=1.52e-06 PS=7.4e-07
mXI0.XI134.MM2 N_XI0.XI134.NET10_XI0.XI134.MM2_d
+ N_XI0.XI134.NET43_XI0.XI134.MM2_g N_VSS_XI0.XI134.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.2375e-13 AS=3.225e-13
+ PD=8.95e-07 PS=1.79e-06
mXI0.XI153.XI0.MM2 N_XI0.G15_XI0.XI153.XI0.MM2_d
+ N_XI0.XI153.NET6_XI0.XI153.XI0.MM2_g N_VSS_XI0.XI153.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI0.XI154.XI0.MM2 N_XI0.G14_XI0.XI154.XI0.MM2_d
+ N_XI0.XI154.NET6_XI0.XI154.XI0.MM2_g N_VSS_XI0.XI154.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI0.XI157.XI0.MM2 N_XI0.G13_XI0.XI157.XI0.MM2_d
+ N_XI0.XI157.NET6_XI0.XI157.XI0.MM2_g N_VSS_XI0.XI157.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI0.XI156.XI0.MM2 N_XI0.G12_XI0.XI156.XI0.MM2_d
+ N_XI0.XI156.NET6_XI0.XI156.XI0.MM2_g N_VSS_XI0.XI156.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI0.XI155.XI0.MM2 N_XI0.G11_XI0.XI155.XI0.MM2_d
+ N_XI0.XI155.NET6_XI0.XI155.XI0.MM2_g N_VSS_XI0.XI155.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI0.XI133.XI0.MM2 N_XI0.G10_XI0.XI133.XI0.MM2_d
+ N_XI0.XI133.NET6_XI0.XI133.XI0.MM2_g N_VSS_XI0.XI133.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI0.XI132.XI0.MM2 N_XI0.G9_XI0.XI132.XI0.MM2_d
+ N_XI0.XI132.NET6_XI0.XI132.XI0.MM2_g N_VSS_XI0.XI132.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI0.XI131.XI0.MM2 N_XI0.G8_XI0.XI131.XI0.MM2_d
+ N_XI0.XI131.NET6_XI0.XI131.XI0.MM2_g N_VSS_XI0.XI131.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI0.XI111.XI0.MM2 N_XI0.G7_XI0.XI111.XI0.MM2_d
+ N_XI0.XI111.NET6_XI0.XI111.XI0.MM2_g N_VSS_XI0.XI111.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI0.XI110.XI0.MM2 N_XI0.G6_XI0.XI110.XI0.MM2_d
+ N_XI0.XI110.NET6_XI0.XI110.XI0.MM2_g N_VSS_XI0.XI110.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI0.XI103.XI0.MM2 N_XI0.G5_XI0.XI103.XI0.MM2_d
+ N_XI0.XI103.NET6_XI0.XI103.XI0.MM2_g N_VSS_XI0.XI103.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI0.XI102.XI0.MM2 N_XI0.G4_XI0.XI102.XI0.MM2_d
+ N_XI0.XI102.NET6_XI0.XI102.XI0.MM2_g N_VSS_XI0.XI102.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI0.XI88.XI0.MM2 N_XI0.G3_XI0.XI88.XI0.MM2_d N_XI0.XI88.NET6_XI0.XI88.XI0.MM2_g
+ N_VSS_XI0.XI88.XI0.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI0.XI82.XI0.MM2 N_XI0.G2_XI0.XI82.XI0.MM2_d N_XI0.XI82.NET6_XI0.XI82.XI0.MM2_g
+ N_VSS_XI0.XI82.XI0.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI0.XI10.XI0.MM2 N_XI0.G1_XI0.XI10.XI0.MM2_d N_XI0.XI10.NET6_XI0.XI10.XI0.MM2_g
+ N_VSS_XI0.XI10.XI0.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI0.XI134.MM7 N_XI0.P16_XI0.XI134.MM7_d N_XI0.XI134.NET39_XI0.XI134.MM7_g
+ N_XI0.XI134.NET10_XI0.XI134.MM7_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=4.75e-13 AS=2.2375e-13 PD=1.9e-06 PS=8.95e-07
mXI0.XI137.XI9.MM2 N_XI0.XI137.NET43_XI0.XI137.XI9.MM2_d
+ N_NET595_XI0.XI137.XI9.MM2_g N_VSS_XI0.XI137.XI9.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI0.XI140.XI9.MM2 N_XI0.XI140.NET43_XI0.XI140.XI9.MM2_d
+ N_NET596_XI0.XI140.XI9.MM2_g N_VSS_XI0.XI140.XI9.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI0.XI149.XI9.MM2 N_XI0.XI149.NET43_XI0.XI149.XI9.MM2_d
+ N_NET597_XI0.XI149.XI9.MM2_g N_VSS_XI0.XI149.XI9.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI0.XI146.XI9.MM2 N_XI0.XI146.NET43_XI0.XI146.XI9.MM2_d
+ N_NET598_XI0.XI146.XI9.MM2_g N_VSS_XI0.XI146.XI9.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI0.XI143.XI9.MM2 N_XI0.XI143.NET43_XI0.XI143.XI9.MM2_d
+ N_NET599_XI0.XI143.XI9.MM2_g N_VSS_XI0.XI143.XI9.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI0.XI128.XI9.MM2 N_XI0.XI128.NET43_XI0.XI128.XI9.MM2_d
+ N_NET600_XI0.XI128.XI9.MM2_g N_VSS_XI0.XI128.XI9.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI0.XI125.XI9.MM2 N_XI0.XI125.NET43_XI0.XI125.XI9.MM2_d
+ N_NET601_XI0.XI125.XI9.MM2_g N_VSS_XI0.XI125.XI9.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI0.XI122.XI9.MM2 N_XI0.XI122.NET43_XI0.XI122.XI9.MM2_d
+ N_NET602_XI0.XI122.XI9.MM2_g N_VSS_XI0.XI122.XI9.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI0.XI114.XI9.MM2 N_XI0.XI114.NET43_XI0.XI114.XI9.MM2_d
+ N_NET603_XI0.XI114.XI9.MM2_g N_VSS_XI0.XI114.XI9.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI0.XI109.XI9.MM2 N_XI0.XI109.NET43_XI0.XI109.XI9.MM2_d
+ N_NET604_XI0.XI109.XI9.MM2_g N_VSS_XI0.XI109.XI9.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI0.XI106.XI9.MM2 N_XI0.XI106.NET43_XI0.XI106.XI9.MM2_d
+ N_NET605_XI0.XI106.XI9.MM2_g N_VSS_XI0.XI106.XI9.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI0.XI101.XI9.MM2 N_XI0.XI101.NET43_XI0.XI101.XI9.MM2_d
+ N_NET606_XI0.XI101.XI9.MM2_g N_VSS_XI0.XI101.XI9.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI0.XI86.XI9.MM2 N_XI0.XI86.NET43_XI0.XI86.XI9.MM2_d
+ N_NET607_XI0.XI86.XI9.MM2_g N_VSS_XI0.XI86.XI9.MM2_s N_VSS_XI10.XI0.XI0.MM2_b
+ N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI0.XI80.XI9.MM2 N_XI0.XI80.NET43_XI0.XI80.XI9.MM2_d
+ N_NET608_XI0.XI80.XI9.MM2_g N_VSS_XI0.XI80.XI9.MM2_s N_VSS_XI10.XI0.XI0.MM2_b
+ N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI0.XI26.XI9.MM2 N_XI0.XI26.NET43_XI0.XI26.XI9.MM2_d
+ N_NET609_XI0.XI26.XI9.MM2_g N_VSS_XI0.XI26.XI9.MM2_s N_VSS_XI10.XI0.XI0.MM2_b
+ N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI0.XI134.MM6 N_XI0.P16_XI0.XI134.MM6_d N_MIN15_XI0.XI134.MM6_g
+ N_XI0.XI134.NET6_XI0.XI134.MM6_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=4.75e-13 AS=1.8125e-13 PD=1.9e-06 PS=7.25e-07
mXI0.XI134.MM0 N_XI0.XI134.NET6_XI0.XI134.MM0_d N_NET594_XI0.XI134.MM0_g
+ N_VSS_XI0.XI134.MM0_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=1.8125e-13 AS=2.575e-13 PD=7.25e-07 PS=1.53e-06
mXI0.XI137.MM2 N_XI0.XI137.NET10_XI0.XI137.MM2_d
+ N_XI0.XI137.NET43_XI0.XI137.MM2_g N_VSS_XI0.XI137.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.2375e-13 AS=3.225e-13
+ PD=8.95e-07 PS=1.79e-06
mXI0.XI140.MM2 N_XI0.XI140.NET10_XI0.XI140.MM2_d
+ N_XI0.XI140.NET43_XI0.XI140.MM2_g N_VSS_XI0.XI140.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.2375e-13 AS=3.225e-13
+ PD=8.95e-07 PS=1.79e-06
mXI0.XI149.MM2 N_XI0.XI149.NET10_XI0.XI149.MM2_d
+ N_XI0.XI149.NET43_XI0.XI149.MM2_g N_VSS_XI0.XI149.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.2375e-13 AS=3.225e-13
+ PD=8.95e-07 PS=1.79e-06
mXI0.XI146.MM2 N_XI0.XI146.NET10_XI0.XI146.MM2_d
+ N_XI0.XI146.NET43_XI0.XI146.MM2_g N_VSS_XI0.XI146.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.2375e-13 AS=3.225e-13
+ PD=8.95e-07 PS=1.79e-06
mXI0.XI143.MM2 N_XI0.XI143.NET10_XI0.XI143.MM2_d
+ N_XI0.XI143.NET43_XI0.XI143.MM2_g N_VSS_XI0.XI143.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.2375e-13 AS=3.225e-13
+ PD=8.95e-07 PS=1.79e-06
mXI0.XI128.MM2 N_XI0.XI128.NET10_XI0.XI128.MM2_d
+ N_XI0.XI128.NET43_XI0.XI128.MM2_g N_VSS_XI0.XI128.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.2375e-13 AS=3.225e-13
+ PD=8.95e-07 PS=1.79e-06
mXI0.XI125.MM2 N_XI0.XI125.NET10_XI0.XI125.MM2_d
+ N_XI0.XI125.NET43_XI0.XI125.MM2_g N_VSS_XI0.XI125.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.2375e-13 AS=3.225e-13
+ PD=8.95e-07 PS=1.79e-06
mXI0.XI122.MM2 N_XI0.XI122.NET10_XI0.XI122.MM2_d
+ N_XI0.XI122.NET43_XI0.XI122.MM2_g N_VSS_XI0.XI122.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.2375e-13 AS=3.225e-13
+ PD=8.95e-07 PS=1.79e-06
mXI0.XI114.MM2 N_XI0.XI114.NET10_XI0.XI114.MM2_d
+ N_XI0.XI114.NET43_XI0.XI114.MM2_g N_VSS_XI0.XI114.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.2375e-13 AS=3.225e-13
+ PD=8.95e-07 PS=1.79e-06
mXI0.XI109.MM2 N_XI0.XI109.NET10_XI0.XI109.MM2_d
+ N_XI0.XI109.NET43_XI0.XI109.MM2_g N_VSS_XI0.XI109.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.2375e-13 AS=3.225e-13
+ PD=8.95e-07 PS=1.79e-06
mXI0.XI106.MM2 N_XI0.XI106.NET10_XI0.XI106.MM2_d
+ N_XI0.XI106.NET43_XI0.XI106.MM2_g N_VSS_XI0.XI106.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.2375e-13 AS=3.225e-13
+ PD=8.95e-07 PS=1.79e-06
mXI0.XI101.MM2 N_XI0.XI101.NET10_XI0.XI101.MM2_d
+ N_XI0.XI101.NET43_XI0.XI101.MM2_g N_VSS_XI0.XI101.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.2375e-13 AS=3.225e-13
+ PD=8.95e-07 PS=1.79e-06
mXI0.XI86.MM2 N_XI0.XI86.NET10_XI0.XI86.MM2_d N_XI0.XI86.NET43_XI0.XI86.MM2_g
+ N_VSS_XI0.XI86.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.2375e-13 AS=3.225e-13 PD=8.95e-07 PS=1.79e-06
mXI0.XI80.MM2 N_XI0.XI80.NET10_XI0.XI80.MM2_d N_XI0.XI80.NET43_XI0.XI80.MM2_g
+ N_VSS_XI0.XI80.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.2375e-13 AS=3.225e-13 PD=8.95e-07 PS=1.79e-06
mXI0.XI26.MM2 N_XI0.XI26.NET10_XI0.XI26.MM2_d N_XI0.XI26.NET43_XI0.XI26.MM2_g
+ N_VSS_XI0.XI26.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.2375e-13 AS=3.225e-13 PD=8.95e-07 PS=1.79e-06
mXI0.XI137.MM7 N_XI0.P15_XI0.XI137.MM7_d N_XI0.XI137.NET39_XI0.XI137.MM7_g
+ N_XI0.XI137.NET10_XI0.XI137.MM7_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=4.75e-13 AS=2.2375e-13 PD=1.9e-06 PS=8.95e-07
mXI0.XI140.MM7 N_XI0.P14_XI0.XI140.MM7_d N_XI0.XI140.NET39_XI0.XI140.MM7_g
+ N_XI0.XI140.NET10_XI0.XI140.MM7_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=4.75e-13 AS=2.2375e-13 PD=1.9e-06 PS=8.95e-07
mXI0.XI149.MM7 N_XI0.P13_XI0.XI149.MM7_d N_XI0.XI149.NET39_XI0.XI149.MM7_g
+ N_XI0.XI149.NET10_XI0.XI149.MM7_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=4.75e-13 AS=2.2375e-13 PD=1.9e-06 PS=8.95e-07
mXI0.XI146.MM7 N_XI0.P12_XI0.XI146.MM7_d N_XI0.XI146.NET39_XI0.XI146.MM7_g
+ N_XI0.XI146.NET10_XI0.XI146.MM7_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=4.75e-13 AS=2.2375e-13 PD=1.9e-06 PS=8.95e-07
mXI0.XI143.MM7 N_XI0.P11_XI0.XI143.MM7_d N_XI0.XI143.NET39_XI0.XI143.MM7_g
+ N_XI0.XI143.NET10_XI0.XI143.MM7_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=4.75e-13 AS=2.2375e-13 PD=1.9e-06 PS=8.95e-07
mXI0.XI128.MM7 N_XI0.P10_XI0.XI128.MM7_d N_XI0.XI128.NET39_XI0.XI128.MM7_g
+ N_XI0.XI128.NET10_XI0.XI128.MM7_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=4.75e-13 AS=2.2375e-13 PD=1.9e-06 PS=8.95e-07
mXI0.XI125.MM7 N_XI0.P9_XI0.XI125.MM7_d N_XI0.XI125.NET39_XI0.XI125.MM7_g
+ N_XI0.XI125.NET10_XI0.XI125.MM7_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=4.75e-13 AS=2.2375e-13 PD=1.9e-06 PS=8.95e-07
mXI0.XI122.MM7 N_XI0.P8_XI0.XI122.MM7_d N_XI0.XI122.NET39_XI0.XI122.MM7_g
+ N_XI0.XI122.NET10_XI0.XI122.MM7_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=4.75e-13 AS=2.2375e-13 PD=1.9e-06 PS=8.95e-07
mXI0.XI114.MM7 N_XI0.P7_XI0.XI114.MM7_d N_XI0.XI114.NET39_XI0.XI114.MM7_g
+ N_XI0.XI114.NET10_XI0.XI114.MM7_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=4.75e-13 AS=2.2375e-13 PD=1.9e-06 PS=8.95e-07
mXI0.XI109.MM7 N_XI0.P6_XI0.XI109.MM7_d N_XI0.XI109.NET39_XI0.XI109.MM7_g
+ N_XI0.XI109.NET10_XI0.XI109.MM7_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=4.75e-13 AS=2.2375e-13 PD=1.9e-06 PS=8.95e-07
mXI0.XI106.MM7 N_XI0.P5_XI0.XI106.MM7_d N_XI0.XI106.NET39_XI0.XI106.MM7_g
+ N_XI0.XI106.NET10_XI0.XI106.MM7_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=4.75e-13 AS=2.2375e-13 PD=1.9e-06 PS=8.95e-07
mXI0.XI101.MM7 N_XI0.P4_XI0.XI101.MM7_d N_XI0.XI101.NET39_XI0.XI101.MM7_g
+ N_XI0.XI101.NET10_XI0.XI101.MM7_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=4.75e-13 AS=2.2375e-13 PD=1.9e-06 PS=8.95e-07
mXI0.XI86.MM7 N_XI0.P3_XI0.XI86.MM7_d N_XI0.XI86.NET39_XI0.XI86.MM7_g
+ N_XI0.XI86.NET10_XI0.XI86.MM7_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=4.75e-13 AS=2.2375e-13 PD=1.9e-06 PS=8.95e-07
mXI0.XI80.MM7 N_XI0.P2_XI0.XI80.MM7_d N_XI0.XI80.NET39_XI0.XI80.MM7_g
+ N_XI0.XI80.NET10_XI0.XI80.MM7_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=4.75e-13 AS=2.2375e-13 PD=1.9e-06 PS=8.95e-07
mXI0.XI26.MM7 N_XI0.P1_XI0.XI26.MM7_d N_XI0.XI26.NET39_XI0.XI26.MM7_g
+ N_XI0.XI26.NET10_XI0.XI26.MM7_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=4.75e-13 AS=2.2375e-13 PD=1.9e-06 PS=8.95e-07
mXI0.XI134.XI4.MM2 N_XI0.XI134.NET39_XI0.XI134.XI4.MM2_d
+ N_MIN15_XI0.XI134.XI4.MM2_g N_VSS_XI0.XI134.XI4.MM2_s N_VSS_XI10.XI0.XI0.MM2_b
+ N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI0.XI137.MM6 N_XI0.P15_XI0.XI137.MM6_d N_MIN14_XI0.XI137.MM6_g
+ N_XI0.XI137.NET6_XI0.XI137.MM6_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=4.75e-13 AS=1.8125e-13 PD=1.9e-06 PS=7.25e-07
mXI0.XI140.MM6 N_XI0.P14_XI0.XI140.MM6_d N_MIN13_XI0.XI140.MM6_g
+ N_XI0.XI140.NET6_XI0.XI140.MM6_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=4.75e-13 AS=1.8125e-13 PD=1.9e-06 PS=7.25e-07
mXI0.XI149.MM6 N_XI0.P13_XI0.XI149.MM6_d N_MIN12_XI0.XI149.MM6_g
+ N_XI0.XI149.NET6_XI0.XI149.MM6_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=4.75e-13 AS=1.8125e-13 PD=1.9e-06 PS=7.25e-07
mXI0.XI146.MM6 N_XI0.P12_XI0.XI146.MM6_d N_MIN11_XI0.XI146.MM6_g
+ N_XI0.XI146.NET6_XI0.XI146.MM6_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=4.75e-13 AS=1.8125e-13 PD=1.9e-06 PS=7.25e-07
mXI0.XI143.MM6 N_XI0.P11_XI0.XI143.MM6_d N_MIN10_XI0.XI143.MM6_g
+ N_XI0.XI143.NET6_XI0.XI143.MM6_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=4.75e-13 AS=1.8125e-13 PD=1.9e-06 PS=7.25e-07
mXI0.XI128.MM6 N_XI0.P10_XI0.XI128.MM6_d N_MIN9_XI0.XI128.MM6_g
+ N_XI0.XI128.NET6_XI0.XI128.MM6_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=4.75e-13 AS=1.8125e-13 PD=1.9e-06 PS=7.25e-07
mXI0.XI125.MM6 N_XI0.P9_XI0.XI125.MM6_d N_MIN8_XI0.XI125.MM6_g
+ N_XI0.XI125.NET6_XI0.XI125.MM6_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=4.75e-13 AS=1.8125e-13 PD=1.9e-06 PS=7.25e-07
mXI0.XI122.MM6 N_XI0.P8_XI0.XI122.MM6_d N_MIN7_XI0.XI122.MM6_g
+ N_XI0.XI122.NET6_XI0.XI122.MM6_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=4.75e-13 AS=1.8125e-13 PD=1.9e-06 PS=7.25e-07
mXI0.XI114.MM6 N_XI0.P7_XI0.XI114.MM6_d N_MIN6_XI0.XI114.MM6_g
+ N_XI0.XI114.NET6_XI0.XI114.MM6_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=4.75e-13 AS=1.8125e-13 PD=1.9e-06 PS=7.25e-07
mXI0.XI109.MM6 N_XI0.P6_XI0.XI109.MM6_d N_MIN5_XI0.XI109.MM6_g
+ N_XI0.XI109.NET6_XI0.XI109.MM6_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=4.75e-13 AS=1.8125e-13 PD=1.9e-06 PS=7.25e-07
mXI0.XI106.MM6 N_XI0.P5_XI0.XI106.MM6_d N_MIN4_XI0.XI106.MM6_g
+ N_XI0.XI106.NET6_XI0.XI106.MM6_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=4.75e-13 AS=1.8125e-13 PD=1.9e-06 PS=7.25e-07
mXI0.XI101.MM6 N_XI0.P4_XI0.XI101.MM6_d N_MIN3_XI0.XI101.MM6_g
+ N_XI0.XI101.NET6_XI0.XI101.MM6_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=4.75e-13 AS=1.8125e-13 PD=1.9e-06 PS=7.25e-07
mXI0.XI86.MM6 N_XI0.P3_XI0.XI86.MM6_d N_MIN2_XI0.XI86.MM6_g
+ N_XI0.XI86.NET6_XI0.XI86.MM6_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=4.75e-13 AS=1.8125e-13 PD=1.9e-06 PS=7.25e-07
mXI0.XI80.MM6 N_XI0.P2_XI0.XI80.MM6_d N_MIN1_XI0.XI80.MM6_g
+ N_XI0.XI80.NET6_XI0.XI80.MM6_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=4.75e-13 AS=1.8125e-13 PD=1.9e-06 PS=7.25e-07
mXI0.XI26.MM6 N_XI0.P1_XI0.XI26.MM6_d N_MIN0_XI0.XI26.MM6_g
+ N_XI0.XI26.NET6_XI0.XI26.MM6_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=4.75e-13 AS=1.8125e-13 PD=1.9e-06 PS=7.25e-07
mXI0.XI137.MM0 N_XI0.XI137.NET6_XI0.XI137.MM0_d N_NET595_XI0.XI137.MM0_g
+ N_VSS_XI0.XI137.MM0_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=1.8125e-13 AS=2.575e-13 PD=7.25e-07 PS=1.53e-06
mXI0.XI140.MM0 N_XI0.XI140.NET6_XI0.XI140.MM0_d N_NET596_XI0.XI140.MM0_g
+ N_VSS_XI0.XI140.MM0_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=1.8125e-13 AS=2.575e-13 PD=7.25e-07 PS=1.53e-06
mXI0.XI149.MM0 N_XI0.XI149.NET6_XI0.XI149.MM0_d N_NET597_XI0.XI149.MM0_g
+ N_VSS_XI0.XI149.MM0_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=1.8125e-13 AS=2.575e-13 PD=7.25e-07 PS=1.53e-06
mXI0.XI146.MM0 N_XI0.XI146.NET6_XI0.XI146.MM0_d N_NET598_XI0.XI146.MM0_g
+ N_VSS_XI0.XI146.MM0_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=1.8125e-13 AS=2.575e-13 PD=7.25e-07 PS=1.53e-06
mXI0.XI143.MM0 N_XI0.XI143.NET6_XI0.XI143.MM0_d N_NET599_XI0.XI143.MM0_g
+ N_VSS_XI0.XI143.MM0_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=1.8125e-13 AS=2.575e-13 PD=7.25e-07 PS=1.53e-06
mXI0.XI128.MM0 N_XI0.XI128.NET6_XI0.XI128.MM0_d N_NET600_XI0.XI128.MM0_g
+ N_VSS_XI0.XI128.MM0_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=1.8125e-13 AS=2.575e-13 PD=7.25e-07 PS=1.53e-06
mXI0.XI125.MM0 N_XI0.XI125.NET6_XI0.XI125.MM0_d N_NET601_XI0.XI125.MM0_g
+ N_VSS_XI0.XI125.MM0_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=1.8125e-13 AS=2.575e-13 PD=7.25e-07 PS=1.53e-06
mXI0.XI122.MM0 N_XI0.XI122.NET6_XI0.XI122.MM0_d N_NET602_XI0.XI122.MM0_g
+ N_VSS_XI0.XI122.MM0_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=1.8125e-13 AS=2.575e-13 PD=7.25e-07 PS=1.53e-06
mXI0.XI114.MM0 N_XI0.XI114.NET6_XI0.XI114.MM0_d N_NET603_XI0.XI114.MM0_g
+ N_VSS_XI0.XI114.MM0_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=1.8125e-13 AS=2.575e-13 PD=7.25e-07 PS=1.53e-06
mXI0.XI109.MM0 N_XI0.XI109.NET6_XI0.XI109.MM0_d N_NET604_XI0.XI109.MM0_g
+ N_VSS_XI0.XI109.MM0_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=1.8125e-13 AS=2.575e-13 PD=7.25e-07 PS=1.53e-06
mXI0.XI106.MM0 N_XI0.XI106.NET6_XI0.XI106.MM0_d N_NET605_XI0.XI106.MM0_g
+ N_VSS_XI0.XI106.MM0_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=1.8125e-13 AS=2.575e-13 PD=7.25e-07 PS=1.53e-06
mXI0.XI101.MM0 N_XI0.XI101.NET6_XI0.XI101.MM0_d N_NET606_XI0.XI101.MM0_g
+ N_VSS_XI0.XI101.MM0_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=1.8125e-13 AS=2.575e-13 PD=7.25e-07 PS=1.53e-06
mXI0.XI86.MM0 N_XI0.XI86.NET6_XI0.XI86.MM0_d N_NET607_XI0.XI86.MM0_g
+ N_VSS_XI0.XI86.MM0_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=1.8125e-13 AS=2.575e-13 PD=7.25e-07 PS=1.53e-06
mXI0.XI80.MM0 N_XI0.XI80.NET6_XI0.XI80.MM0_d N_NET608_XI0.XI80.MM0_g
+ N_VSS_XI0.XI80.MM0_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=1.8125e-13 AS=2.575e-13 PD=7.25e-07 PS=1.53e-06
mXI0.XI26.MM0 N_XI0.XI26.NET6_XI0.XI26.MM0_d N_NET609_XI0.XI26.MM0_g
+ N_VSS_XI0.XI26.MM0_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=1.8125e-13 AS=2.575e-13 PD=7.25e-07 PS=1.53e-06
mXI6.MM2 N_NET0859_XI6.MM2_d N_NET0858_XI6.MM2_g N_VSS_XI6.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=3e-06 AD=1.47e-12 AS=1.47e-12
+ PD=3.98e-06 PS=3.98e-06
mXI0.XI182.XI9.MM2 N_XI0.XI182.NET43_XI0.XI182.XI9.MM2_d
+ N_XI0.P16_XI0.XI182.XI9.MM2_g N_VSS_XI0.XI182.XI9.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI0.XI137.XI4.MM2 N_XI0.XI137.NET39_XI0.XI137.XI4.MM2_d
+ N_MIN14_XI0.XI137.XI4.MM2_g N_VSS_XI0.XI137.XI4.MM2_s N_VSS_XI10.XI0.XI0.MM2_b
+ N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI0.XI140.XI4.MM2 N_XI0.XI140.NET39_XI0.XI140.XI4.MM2_d
+ N_MIN13_XI0.XI140.XI4.MM2_g N_VSS_XI0.XI140.XI4.MM2_s N_VSS_XI10.XI0.XI0.MM2_b
+ N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI0.XI149.XI4.MM2 N_XI0.XI149.NET39_XI0.XI149.XI4.MM2_d
+ N_MIN12_XI0.XI149.XI4.MM2_g N_VSS_XI0.XI149.XI4.MM2_s N_VSS_XI10.XI0.XI0.MM2_b
+ N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI0.XI146.XI4.MM2 N_XI0.XI146.NET39_XI0.XI146.XI4.MM2_d
+ N_MIN11_XI0.XI146.XI4.MM2_g N_VSS_XI0.XI146.XI4.MM2_s N_VSS_XI10.XI0.XI0.MM2_b
+ N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI0.XI143.XI4.MM2 N_XI0.XI143.NET39_XI0.XI143.XI4.MM2_d
+ N_MIN10_XI0.XI143.XI4.MM2_g N_VSS_XI0.XI143.XI4.MM2_s N_VSS_XI10.XI0.XI0.MM2_b
+ N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI0.XI128.XI4.MM2 N_XI0.XI128.NET39_XI0.XI128.XI4.MM2_d
+ N_MIN9_XI0.XI128.XI4.MM2_g N_VSS_XI0.XI128.XI4.MM2_s N_VSS_XI10.XI0.XI0.MM2_b
+ N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI0.XI125.XI4.MM2 N_XI0.XI125.NET39_XI0.XI125.XI4.MM2_d
+ N_MIN8_XI0.XI125.XI4.MM2_g N_VSS_XI0.XI125.XI4.MM2_s N_VSS_XI10.XI0.XI0.MM2_b
+ N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI0.XI122.XI4.MM2 N_XI0.XI122.NET39_XI0.XI122.XI4.MM2_d
+ N_MIN7_XI0.XI122.XI4.MM2_g N_VSS_XI0.XI122.XI4.MM2_s N_VSS_XI10.XI0.XI0.MM2_b
+ N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI0.XI114.XI4.MM2 N_XI0.XI114.NET39_XI0.XI114.XI4.MM2_d
+ N_MIN6_XI0.XI114.XI4.MM2_g N_VSS_XI0.XI114.XI4.MM2_s N_VSS_XI10.XI0.XI0.MM2_b
+ N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI0.XI109.XI4.MM2 N_XI0.XI109.NET39_XI0.XI109.XI4.MM2_d
+ N_MIN5_XI0.XI109.XI4.MM2_g N_VSS_XI0.XI109.XI4.MM2_s N_VSS_XI10.XI0.XI0.MM2_b
+ N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI0.XI106.XI4.MM2 N_XI0.XI106.NET39_XI0.XI106.XI4.MM2_d
+ N_MIN4_XI0.XI106.XI4.MM2_g N_VSS_XI0.XI106.XI4.MM2_s N_VSS_XI10.XI0.XI0.MM2_b
+ N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI0.XI101.XI4.MM2 N_XI0.XI101.NET39_XI0.XI101.XI4.MM2_d
+ N_MIN3_XI0.XI101.XI4.MM2_g N_VSS_XI0.XI101.XI4.MM2_s N_VSS_XI10.XI0.XI0.MM2_b
+ N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI0.XI86.XI4.MM2 N_XI0.XI86.NET39_XI0.XI86.XI4.MM2_d N_MIN2_XI0.XI86.XI4.MM2_g
+ N_VSS_XI0.XI86.XI4.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI0.XI80.XI4.MM2 N_XI0.XI80.NET39_XI0.XI80.XI4.MM2_d N_MIN1_XI0.XI80.XI4.MM2_g
+ N_VSS_XI0.XI80.XI4.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI0.XI26.XI4.MM2 N_XI0.XI26.NET39_XI0.XI26.XI4.MM2_d N_MIN0_XI0.XI26.XI4.MM2_g
+ N_VSS_XI0.XI26.XI4.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI0.XI182.MM2 N_XI0.XI182.NET10_XI0.XI182.MM2_d
+ N_XI0.XI182.NET43_XI0.XI182.MM2_g N_VSS_XI0.XI182.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.2375e-13 AS=3.225e-13
+ PD=8.95e-07 PS=1.79e-06
mXI0.XI168.XI1.XI1.MM0 N_XI0.XI168.XI1.XI1.NET036_XI0.XI168.XI1.XI1.MM0_d
+ N_XI0.NET288_XI0.XI168.XI1.XI1.MM0_g N_VSS_XI0.XI168.XI1.XI1.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.85e-13 AS=2.45e-13
+ PD=7.4e-07 PS=1.48e-06
mXI0.XI167.XI1.XI1.MM0 N_XI0.XI167.XI1.XI1.NET036_XI0.XI167.XI1.XI1.MM0_d
+ N_XI0.NET282_XI0.XI167.XI1.XI1.MM0_g N_VSS_XI0.XI167.XI1.XI1.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.85e-13 AS=2.45e-13
+ PD=7.4e-07 PS=1.48e-06
mXI0.XI166.XI1.XI1.MM0 N_XI0.XI166.XI1.XI1.NET036_XI0.XI166.XI1.XI1.MM0_d
+ N_XI0.NET276_XI0.XI166.XI1.XI1.MM0_g N_VSS_XI0.XI166.XI1.XI1.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.85e-13 AS=2.45e-13
+ PD=7.4e-07 PS=1.48e-06
mXI0.XI165.XI1.XI1.MM0 N_XI0.XI165.XI1.XI1.NET036_XI0.XI165.XI1.XI1.MM0_d
+ N_XI0.NET270_XI0.XI165.XI1.XI1.MM0_g N_VSS_XI0.XI165.XI1.XI1.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.85e-13 AS=2.45e-13
+ PD=7.4e-07 PS=1.48e-06
mXI0.XI159.XI1.XI1.MM0 N_XI0.XI159.XI1.XI1.NET036_XI0.XI159.XI1.XI1.MM0_d
+ N_XI0.NET246_XI0.XI159.XI1.XI1.MM0_g N_VSS_XI0.XI159.XI1.XI1.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.85e-13 AS=2.45e-13
+ PD=7.4e-07 PS=1.48e-06
mXI0.XI160.XI1.XI1.MM0 N_XI0.XI160.XI1.XI1.NET036_XI0.XI160.XI1.XI1.MM0_d
+ N_XI0.NET252_XI0.XI160.XI1.XI1.MM0_g N_VSS_XI0.XI160.XI1.XI1.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.85e-13 AS=2.45e-13
+ PD=7.4e-07 PS=1.48e-06
mXI0.XI161.XI1.XI1.MM0 N_XI0.XI161.XI1.XI1.NET036_XI0.XI161.XI1.XI1.MM0_d
+ N_XI0.NET258_XI0.XI161.XI1.XI1.MM0_g N_VSS_XI0.XI161.XI1.XI1.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.85e-13 AS=2.45e-13
+ PD=7.4e-07 PS=1.48e-06
mXI0.XI162.XI1.XI1.MM0 N_XI0.XI162.XI1.XI1.NET036_XI0.XI162.XI1.XI1.MM0_d
+ N_XI0.NET264_XI0.XI162.XI1.XI1.MM0_g N_VSS_XI0.XI162.XI1.XI1.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.85e-13 AS=2.45e-13
+ PD=7.4e-07 PS=1.48e-06
mXI0.XI121.XI1.XI1.MM0 N_XI0.XI121.XI1.XI1.NET036_XI0.XI121.XI1.XI1.MM0_d
+ N_XI0.NET204_XI0.XI121.XI1.XI1.MM0_g N_VSS_XI0.XI121.XI1.XI1.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.85e-13 AS=2.45e-13
+ PD=7.4e-07 PS=1.48e-06
mXI0.XI120.XI1.XI1.MM0 N_XI0.XI120.XI1.XI1.NET036_XI0.XI120.XI1.XI1.MM0_d
+ N_XI0.NET210_XI0.XI120.XI1.XI1.MM0_g N_VSS_XI0.XI120.XI1.XI1.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.85e-13 AS=2.45e-13
+ PD=7.4e-07 PS=1.48e-06
mXI0.XI119.XI1.XI1.MM0 N_XI0.XI119.XI1.XI1.NET036_XI0.XI119.XI1.XI1.MM0_d
+ N_XI0.NET216_XI0.XI119.XI1.XI1.MM0_g N_VSS_XI0.XI119.XI1.XI1.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.85e-13 AS=2.45e-13
+ PD=7.4e-07 PS=1.48e-06
mXI0.XI118.XI1.XI1.MM0 N_XI0.XI118.XI1.XI1.NET036_XI0.XI118.XI1.XI1.MM0_d
+ N_XI0.NET222_XI0.XI118.XI1.XI1.MM0_g N_VSS_XI0.XI118.XI1.XI1.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.85e-13 AS=2.45e-13
+ PD=7.4e-07 PS=1.48e-06
mXI0.XI91.XI1.XI1.MM0 N_XI0.XI91.XI1.XI1.NET036_XI0.XI91.XI1.XI1.MM0_d
+ N_XI0.NET228_XI0.XI91.XI1.XI1.MM0_g N_VSS_XI0.XI91.XI1.XI1.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.85e-13 AS=2.45e-13
+ PD=7.4e-07 PS=1.48e-06
mXI0.XI90.XI1.XI1.MM0 N_XI0.XI90.XI1.XI1.NET036_XI0.XI90.XI1.XI1.MM0_d
+ N_XI0.NET240_XI0.XI90.XI1.XI1.MM0_g N_VSS_XI0.XI90.XI1.XI1.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.85e-13 AS=2.45e-13
+ PD=7.4e-07 PS=1.48e-06
mXI0.XI89.XI1.XI1.MM0 N_XI0.XI89.XI1.XI1.NET036_XI0.XI89.XI1.XI1.MM0_d
+ N_CIN2_XI0.XI89.XI1.XI1.MM0_g N_VSS_XI0.XI89.XI1.XI1.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.85e-13 AS=2.45e-13
+ PD=7.4e-07 PS=1.48e-06
mXI0.XI182.MM7 N_NET141_XI0.XI182.MM7_d N_XI0.XI182.NET39_XI0.XI182.MM7_g
+ N_XI0.XI182.NET10_XI0.XI182.MM7_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=4.75e-13 AS=2.2375e-13 PD=1.9e-06 PS=8.95e-07
mXI0.XI168.XI1.XI1.MM2 N_XI0.XI168.XI1.NET6_XI0.XI168.XI1.XI1.MM2_d
+ N_XI0.P15_XI0.XI168.XI1.XI1.MM2_g
+ N_XI0.XI168.XI1.XI1.NET036_XI0.XI168.XI1.XI1.MM2_s N_VSS_XI10.XI0.XI0.MM2_b
+ N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=1.85e-13 PD=1.52e-06 PS=7.4e-07
mXI0.XI167.XI1.XI1.MM2 N_XI0.XI167.XI1.NET6_XI0.XI167.XI1.XI1.MM2_d
+ N_XI0.P14_XI0.XI167.XI1.XI1.MM2_g
+ N_XI0.XI167.XI1.XI1.NET036_XI0.XI167.XI1.XI1.MM2_s N_VSS_XI10.XI0.XI0.MM2_b
+ N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=1.85e-13 PD=1.52e-06 PS=7.4e-07
mXI0.XI166.XI1.XI1.MM2 N_XI0.XI166.XI1.NET6_XI0.XI166.XI1.XI1.MM2_d
+ N_XI0.P13_XI0.XI166.XI1.XI1.MM2_g
+ N_XI0.XI166.XI1.XI1.NET036_XI0.XI166.XI1.XI1.MM2_s N_VSS_XI10.XI0.XI0.MM2_b
+ N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=1.85e-13 PD=1.52e-06 PS=7.4e-07
mXI0.XI165.XI1.XI1.MM2 N_XI0.XI165.XI1.NET6_XI0.XI165.XI1.XI1.MM2_d
+ N_XI0.P12_XI0.XI165.XI1.XI1.MM2_g
+ N_XI0.XI165.XI1.XI1.NET036_XI0.XI165.XI1.XI1.MM2_s N_VSS_XI10.XI0.XI0.MM2_b
+ N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=1.85e-13 PD=1.52e-06 PS=7.4e-07
mXI0.XI159.XI1.XI1.MM2 N_XI0.XI159.XI1.NET6_XI0.XI159.XI1.XI1.MM2_d
+ N_XI0.P11_XI0.XI159.XI1.XI1.MM2_g
+ N_XI0.XI159.XI1.XI1.NET036_XI0.XI159.XI1.XI1.MM2_s N_VSS_XI10.XI0.XI0.MM2_b
+ N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=1.85e-13 PD=1.52e-06 PS=7.4e-07
mXI0.XI160.XI1.XI1.MM2 N_XI0.XI160.XI1.NET6_XI0.XI160.XI1.XI1.MM2_d
+ N_XI0.P10_XI0.XI160.XI1.XI1.MM2_g
+ N_XI0.XI160.XI1.XI1.NET036_XI0.XI160.XI1.XI1.MM2_s N_VSS_XI10.XI0.XI0.MM2_b
+ N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=1.85e-13 PD=1.52e-06 PS=7.4e-07
mXI0.XI161.XI1.XI1.MM2 N_XI0.XI161.XI1.NET6_XI0.XI161.XI1.XI1.MM2_d
+ N_XI0.P9_XI0.XI161.XI1.XI1.MM2_g
+ N_XI0.XI161.XI1.XI1.NET036_XI0.XI161.XI1.XI1.MM2_s N_VSS_XI10.XI0.XI0.MM2_b
+ N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=1.85e-13 PD=1.52e-06 PS=7.4e-07
mXI0.XI162.XI1.XI1.MM2 N_XI0.XI162.XI1.NET6_XI0.XI162.XI1.XI1.MM2_d
+ N_XI0.P8_XI0.XI162.XI1.XI1.MM2_g
+ N_XI0.XI162.XI1.XI1.NET036_XI0.XI162.XI1.XI1.MM2_s N_VSS_XI10.XI0.XI0.MM2_b
+ N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=1.85e-13 PD=1.52e-06 PS=7.4e-07
mXI0.XI121.XI1.XI1.MM2 N_XI0.XI121.XI1.NET6_XI0.XI121.XI1.XI1.MM2_d
+ N_XI0.P7_XI0.XI121.XI1.XI1.MM2_g
+ N_XI0.XI121.XI1.XI1.NET036_XI0.XI121.XI1.XI1.MM2_s N_VSS_XI10.XI0.XI0.MM2_b
+ N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=1.85e-13 PD=1.52e-06 PS=7.4e-07
mXI0.XI120.XI1.XI1.MM2 N_XI0.XI120.XI1.NET6_XI0.XI120.XI1.XI1.MM2_d
+ N_XI0.P6_XI0.XI120.XI1.XI1.MM2_g
+ N_XI0.XI120.XI1.XI1.NET036_XI0.XI120.XI1.XI1.MM2_s N_VSS_XI10.XI0.XI0.MM2_b
+ N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=1.85e-13 PD=1.52e-06 PS=7.4e-07
mXI0.XI119.XI1.XI1.MM2 N_XI0.XI119.XI1.NET6_XI0.XI119.XI1.XI1.MM2_d
+ N_XI0.P5_XI0.XI119.XI1.XI1.MM2_g
+ N_XI0.XI119.XI1.XI1.NET036_XI0.XI119.XI1.XI1.MM2_s N_VSS_XI10.XI0.XI0.MM2_b
+ N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=1.85e-13 PD=1.52e-06 PS=7.4e-07
mXI0.XI118.XI1.XI1.MM2 N_XI0.XI118.XI1.NET6_XI0.XI118.XI1.XI1.MM2_d
+ N_XI0.P4_XI0.XI118.XI1.XI1.MM2_g
+ N_XI0.XI118.XI1.XI1.NET036_XI0.XI118.XI1.XI1.MM2_s N_VSS_XI10.XI0.XI0.MM2_b
+ N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=1.85e-13 PD=1.52e-06 PS=7.4e-07
mXI0.XI91.XI1.XI1.MM2 N_XI0.XI91.XI1.NET6_XI0.XI91.XI1.XI1.MM2_d
+ N_XI0.P3_XI0.XI91.XI1.XI1.MM2_g
+ N_XI0.XI91.XI1.XI1.NET036_XI0.XI91.XI1.XI1.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18
+ L=1.8e-07 W=5e-07 AD=2.55e-13 AS=1.85e-13 PD=1.52e-06 PS=7.4e-07
mXI0.XI90.XI1.XI1.MM2 N_XI0.XI90.XI1.NET6_XI0.XI90.XI1.XI1.MM2_d
+ N_XI0.P2_XI0.XI90.XI1.XI1.MM2_g
+ N_XI0.XI90.XI1.XI1.NET036_XI0.XI90.XI1.XI1.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18
+ L=1.8e-07 W=5e-07 AD=2.55e-13 AS=1.85e-13 PD=1.52e-06 PS=7.4e-07
mXI0.XI89.XI1.XI1.MM2 N_XI0.XI89.XI1.NET6_XI0.XI89.XI1.XI1.MM2_d
+ N_XI0.P1_XI0.XI89.XI1.XI1.MM2_g
+ N_XI0.XI89.XI1.XI1.NET036_XI0.XI89.XI1.XI1.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18
+ L=1.8e-07 W=5e-07 AD=2.55e-13 AS=1.85e-13 PD=1.52e-06 PS=7.4e-07
mXI0.XI182.MM6 N_NET141_XI0.XI182.MM6_d N_XI0.NET198_XI0.XI182.MM6_g
+ N_XI0.XI182.NET6_XI0.XI182.MM6_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=4.75e-13 AS=1.8125e-13 PD=1.9e-06 PS=7.25e-07
mXI0.XI168.XI1.XI0.MM2 N_XI0.XI168.NET13_XI0.XI168.XI1.XI0.MM2_d
+ N_XI0.XI168.XI1.NET6_XI0.XI168.XI1.XI0.MM2_g N_VSS_XI0.XI168.XI1.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI0.XI167.XI1.XI0.MM2 N_XI0.XI167.NET13_XI0.XI167.XI1.XI0.MM2_d
+ N_XI0.XI167.XI1.NET6_XI0.XI167.XI1.XI0.MM2_g N_VSS_XI0.XI167.XI1.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI0.XI166.XI1.XI0.MM2 N_XI0.XI166.NET13_XI0.XI166.XI1.XI0.MM2_d
+ N_XI0.XI166.XI1.NET6_XI0.XI166.XI1.XI0.MM2_g N_VSS_XI0.XI166.XI1.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI0.XI165.XI1.XI0.MM2 N_XI0.XI165.NET13_XI0.XI165.XI1.XI0.MM2_d
+ N_XI0.XI165.XI1.NET6_XI0.XI165.XI1.XI0.MM2_g N_VSS_XI0.XI165.XI1.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI0.XI159.XI1.XI0.MM2 N_XI0.XI159.NET13_XI0.XI159.XI1.XI0.MM2_d
+ N_XI0.XI159.XI1.NET6_XI0.XI159.XI1.XI0.MM2_g N_VSS_XI0.XI159.XI1.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI0.XI160.XI1.XI0.MM2 N_XI0.XI160.NET13_XI0.XI160.XI1.XI0.MM2_d
+ N_XI0.XI160.XI1.NET6_XI0.XI160.XI1.XI0.MM2_g N_VSS_XI0.XI160.XI1.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI0.XI161.XI1.XI0.MM2 N_XI0.XI161.NET13_XI0.XI161.XI1.XI0.MM2_d
+ N_XI0.XI161.XI1.NET6_XI0.XI161.XI1.XI0.MM2_g N_VSS_XI0.XI161.XI1.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI0.XI162.XI1.XI0.MM2 N_XI0.XI162.NET13_XI0.XI162.XI1.XI0.MM2_d
+ N_XI0.XI162.XI1.NET6_XI0.XI162.XI1.XI0.MM2_g N_VSS_XI0.XI162.XI1.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI0.XI121.XI1.XI0.MM2 N_XI0.XI121.NET13_XI0.XI121.XI1.XI0.MM2_d
+ N_XI0.XI121.XI1.NET6_XI0.XI121.XI1.XI0.MM2_g N_VSS_XI0.XI121.XI1.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI0.XI120.XI1.XI0.MM2 N_XI0.XI120.NET13_XI0.XI120.XI1.XI0.MM2_d
+ N_XI0.XI120.XI1.NET6_XI0.XI120.XI1.XI0.MM2_g N_VSS_XI0.XI120.XI1.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI0.XI119.XI1.XI0.MM2 N_XI0.XI119.NET13_XI0.XI119.XI1.XI0.MM2_d
+ N_XI0.XI119.XI1.NET6_XI0.XI119.XI1.XI0.MM2_g N_VSS_XI0.XI119.XI1.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI0.XI118.XI1.XI0.MM2 N_XI0.XI118.NET13_XI0.XI118.XI1.XI0.MM2_d
+ N_XI0.XI118.XI1.NET6_XI0.XI118.XI1.XI0.MM2_g N_VSS_XI0.XI118.XI1.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI0.XI91.XI1.XI0.MM2 N_XI0.XI91.NET13_XI0.XI91.XI1.XI0.MM2_d
+ N_XI0.XI91.XI1.NET6_XI0.XI91.XI1.XI0.MM2_g N_VSS_XI0.XI91.XI1.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI0.XI90.XI1.XI0.MM2 N_XI0.XI90.NET13_XI0.XI90.XI1.XI0.MM2_d
+ N_XI0.XI90.XI1.NET6_XI0.XI90.XI1.XI0.MM2_g N_VSS_XI0.XI90.XI1.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI0.XI89.XI1.XI0.MM2 N_XI0.XI89.NET13_XI0.XI89.XI1.XI0.MM2_d
+ N_XI0.XI89.XI1.NET6_XI0.XI89.XI1.XI0.MM2_g N_VSS_XI0.XI89.XI1.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI0.XI182.MM0 N_XI0.XI182.NET6_XI0.XI182.MM0_d N_XI0.P16_XI0.XI182.MM0_g
+ N_VSS_XI0.XI182.MM0_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=1.8125e-13 AS=2.575e-13 PD=7.25e-07 PS=1.53e-06
mXI0.XI168.XI0.XI0.MM0 N_XI0.XI168.XI0.NET12_XI0.XI168.XI0.XI0.MM0_d
+ N_XI0.XI168.NET13_XI0.XI168.XI0.XI0.MM0_g N_VSS_XI0.XI168.XI0.XI0.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.375e-13 AS=2.45e-13
+ PD=5.5e-07 PS=1.48e-06
mXI0.XI167.XI0.XI0.MM0 N_XI0.XI167.XI0.NET12_XI0.XI167.XI0.XI0.MM0_d
+ N_XI0.XI167.NET13_XI0.XI167.XI0.XI0.MM0_g N_VSS_XI0.XI167.XI0.XI0.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.375e-13 AS=2.45e-13
+ PD=5.5e-07 PS=1.48e-06
mXI0.XI166.XI0.XI0.MM0 N_XI0.XI166.XI0.NET12_XI0.XI166.XI0.XI0.MM0_d
+ N_XI0.XI166.NET13_XI0.XI166.XI0.XI0.MM0_g N_VSS_XI0.XI166.XI0.XI0.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.375e-13 AS=2.45e-13
+ PD=5.5e-07 PS=1.48e-06
mXI0.XI165.XI0.XI0.MM0 N_XI0.XI165.XI0.NET12_XI0.XI165.XI0.XI0.MM0_d
+ N_XI0.XI165.NET13_XI0.XI165.XI0.XI0.MM0_g N_VSS_XI0.XI165.XI0.XI0.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.375e-13 AS=2.45e-13
+ PD=5.5e-07 PS=1.48e-06
mXI0.XI159.XI0.XI0.MM0 N_XI0.XI159.XI0.NET12_XI0.XI159.XI0.XI0.MM0_d
+ N_XI0.XI159.NET13_XI0.XI159.XI0.XI0.MM0_g N_VSS_XI0.XI159.XI0.XI0.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.375e-13 AS=2.45e-13
+ PD=5.5e-07 PS=1.48e-06
mXI0.XI160.XI0.XI0.MM0 N_XI0.XI160.XI0.NET12_XI0.XI160.XI0.XI0.MM0_d
+ N_XI0.XI160.NET13_XI0.XI160.XI0.XI0.MM0_g N_VSS_XI0.XI160.XI0.XI0.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.375e-13 AS=2.45e-13
+ PD=5.5e-07 PS=1.48e-06
mXI0.XI161.XI0.XI0.MM0 N_XI0.XI161.XI0.NET12_XI0.XI161.XI0.XI0.MM0_d
+ N_XI0.XI161.NET13_XI0.XI161.XI0.XI0.MM0_g N_VSS_XI0.XI161.XI0.XI0.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.375e-13 AS=2.45e-13
+ PD=5.5e-07 PS=1.48e-06
mXI0.XI162.XI0.XI0.MM0 N_XI0.XI162.XI0.NET12_XI0.XI162.XI0.XI0.MM0_d
+ N_XI0.XI162.NET13_XI0.XI162.XI0.XI0.MM0_g N_VSS_XI0.XI162.XI0.XI0.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.375e-13 AS=2.45e-13
+ PD=5.5e-07 PS=1.48e-06
mXI0.XI121.XI0.XI0.MM0 N_XI0.XI121.XI0.NET12_XI0.XI121.XI0.XI0.MM0_d
+ N_XI0.XI121.NET13_XI0.XI121.XI0.XI0.MM0_g N_VSS_XI0.XI121.XI0.XI0.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.375e-13 AS=2.45e-13
+ PD=5.5e-07 PS=1.48e-06
mXI0.XI120.XI0.XI0.MM0 N_XI0.XI120.XI0.NET12_XI0.XI120.XI0.XI0.MM0_d
+ N_XI0.XI120.NET13_XI0.XI120.XI0.XI0.MM0_g N_VSS_XI0.XI120.XI0.XI0.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.375e-13 AS=2.45e-13
+ PD=5.5e-07 PS=1.48e-06
mXI0.XI119.XI0.XI0.MM0 N_XI0.XI119.XI0.NET12_XI0.XI119.XI0.XI0.MM0_d
+ N_XI0.XI119.NET13_XI0.XI119.XI0.XI0.MM0_g N_VSS_XI0.XI119.XI0.XI0.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.375e-13 AS=2.45e-13
+ PD=5.5e-07 PS=1.48e-06
mXI0.XI118.XI0.XI0.MM0 N_XI0.XI118.XI0.NET12_XI0.XI118.XI0.XI0.MM0_d
+ N_XI0.XI118.NET13_XI0.XI118.XI0.XI0.MM0_g N_VSS_XI0.XI118.XI0.XI0.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.375e-13 AS=2.45e-13
+ PD=5.5e-07 PS=1.48e-06
mXI0.XI91.XI0.XI0.MM0 N_XI0.XI91.XI0.NET12_XI0.XI91.XI0.XI0.MM0_d
+ N_XI0.XI91.NET13_XI0.XI91.XI0.XI0.MM0_g N_VSS_XI0.XI91.XI0.XI0.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.375e-13 AS=2.45e-13
+ PD=5.5e-07 PS=1.48e-06
mXI0.XI90.XI0.XI0.MM0 N_XI0.XI90.XI0.NET12_XI0.XI90.XI0.XI0.MM0_d
+ N_XI0.XI90.NET13_XI0.XI90.XI0.XI0.MM0_g N_VSS_XI0.XI90.XI0.XI0.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.375e-13 AS=2.45e-13
+ PD=5.5e-07 PS=1.48e-06
mXI0.XI89.XI0.XI0.MM0 N_XI0.XI89.XI0.NET12_XI0.XI89.XI0.XI0.MM0_d
+ N_XI0.XI89.NET13_XI0.XI89.XI0.XI0.MM0_g N_VSS_XI0.XI89.XI0.XI0.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.375e-13 AS=2.45e-13
+ PD=5.5e-07 PS=1.48e-06
mXI0.XI182.XI4.MM2 N_XI0.XI182.NET39_XI0.XI182.XI4.MM2_d
+ N_XI0.NET198_XI0.XI182.XI4.MM2_g N_VSS_XI0.XI182.XI4.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI2.MM2 N_NET0858_XI2.MM2_d N_NET141_XI2.MM2_g N_VSS_XI2.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI0.XI168.XI0.XI0.MM2 N_XI0.XI168.XI0.NET12_XI0.XI168.XI0.XI0.MM2_d
+ N_XI0.G15_XI0.XI168.XI0.XI0.MM2_g N_VSS_XI0.XI168.XI0.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.375e-13 AS=2.55e-13
+ PD=5.5e-07 PS=1.52e-06
mXI0.XI167.XI0.XI0.MM2 N_XI0.XI167.XI0.NET12_XI0.XI167.XI0.XI0.MM2_d
+ N_XI0.G14_XI0.XI167.XI0.XI0.MM2_g N_VSS_XI0.XI167.XI0.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.375e-13 AS=2.55e-13
+ PD=5.5e-07 PS=1.52e-06
mXI0.XI166.XI0.XI0.MM2 N_XI0.XI166.XI0.NET12_XI0.XI166.XI0.XI0.MM2_d
+ N_XI0.G13_XI0.XI166.XI0.XI0.MM2_g N_VSS_XI0.XI166.XI0.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.375e-13 AS=2.55e-13
+ PD=5.5e-07 PS=1.52e-06
mXI0.XI165.XI0.XI0.MM2 N_XI0.XI165.XI0.NET12_XI0.XI165.XI0.XI0.MM2_d
+ N_XI0.G12_XI0.XI165.XI0.XI0.MM2_g N_VSS_XI0.XI165.XI0.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.375e-13 AS=2.55e-13
+ PD=5.5e-07 PS=1.52e-06
mXI0.XI159.XI0.XI0.MM2 N_XI0.XI159.XI0.NET12_XI0.XI159.XI0.XI0.MM2_d
+ N_XI0.G11_XI0.XI159.XI0.XI0.MM2_g N_VSS_XI0.XI159.XI0.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.375e-13 AS=2.55e-13
+ PD=5.5e-07 PS=1.52e-06
mXI0.XI160.XI0.XI0.MM2 N_XI0.XI160.XI0.NET12_XI0.XI160.XI0.XI0.MM2_d
+ N_XI0.G10_XI0.XI160.XI0.XI0.MM2_g N_VSS_XI0.XI160.XI0.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.375e-13 AS=2.55e-13
+ PD=5.5e-07 PS=1.52e-06
mXI0.XI161.XI0.XI0.MM2 N_XI0.XI161.XI0.NET12_XI0.XI161.XI0.XI0.MM2_d
+ N_XI0.G9_XI0.XI161.XI0.XI0.MM2_g N_VSS_XI0.XI161.XI0.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.375e-13 AS=2.55e-13
+ PD=5.5e-07 PS=1.52e-06
mXI0.XI162.XI0.XI0.MM2 N_XI0.XI162.XI0.NET12_XI0.XI162.XI0.XI0.MM2_d
+ N_XI0.G8_XI0.XI162.XI0.XI0.MM2_g N_VSS_XI0.XI162.XI0.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.375e-13 AS=2.55e-13
+ PD=5.5e-07 PS=1.52e-06
mXI0.XI121.XI0.XI0.MM2 N_XI0.XI121.XI0.NET12_XI0.XI121.XI0.XI0.MM2_d
+ N_XI0.G7_XI0.XI121.XI0.XI0.MM2_g N_VSS_XI0.XI121.XI0.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.375e-13 AS=2.55e-13
+ PD=5.5e-07 PS=1.52e-06
mXI0.XI120.XI0.XI0.MM2 N_XI0.XI120.XI0.NET12_XI0.XI120.XI0.XI0.MM2_d
+ N_XI0.G6_XI0.XI120.XI0.XI0.MM2_g N_VSS_XI0.XI120.XI0.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.375e-13 AS=2.55e-13
+ PD=5.5e-07 PS=1.52e-06
mXI0.XI119.XI0.XI0.MM2 N_XI0.XI119.XI0.NET12_XI0.XI119.XI0.XI0.MM2_d
+ N_XI0.G5_XI0.XI119.XI0.XI0.MM2_g N_VSS_XI0.XI119.XI0.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.375e-13 AS=2.55e-13
+ PD=5.5e-07 PS=1.52e-06
mXI0.XI118.XI0.XI0.MM2 N_XI0.XI118.XI0.NET12_XI0.XI118.XI0.XI0.MM2_d
+ N_XI0.G4_XI0.XI118.XI0.XI0.MM2_g N_VSS_XI0.XI118.XI0.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.375e-13 AS=2.55e-13
+ PD=5.5e-07 PS=1.52e-06
mXI0.XI91.XI0.XI0.MM2 N_XI0.XI91.XI0.NET12_XI0.XI91.XI0.XI0.MM2_d
+ N_XI0.G3_XI0.XI91.XI0.XI0.MM2_g N_VSS_XI0.XI91.XI0.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.375e-13 AS=2.55e-13
+ PD=5.5e-07 PS=1.52e-06
mXI0.XI90.XI0.XI0.MM2 N_XI0.XI90.XI0.NET12_XI0.XI90.XI0.XI0.MM2_d
+ N_XI0.G2_XI0.XI90.XI0.XI0.MM2_g N_VSS_XI0.XI90.XI0.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.375e-13 AS=2.55e-13
+ PD=5.5e-07 PS=1.52e-06
mXI0.XI89.XI0.XI0.MM2 N_XI0.XI89.XI0.NET12_XI0.XI89.XI0.XI0.MM2_d
+ N_XI0.G1_XI0.XI89.XI0.XI0.MM2_g N_VSS_XI0.XI89.XI0.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.375e-13 AS=2.55e-13
+ PD=5.5e-07 PS=1.52e-06
mXI0.XI168.XI0.XI1.MM2 N_XI0.NET198_XI0.XI168.XI0.XI1.MM2_d
+ N_XI0.XI168.XI0.NET12_XI0.XI168.XI0.XI1.MM2_g N_VSS_XI0.XI168.XI0.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI0.XI167.XI0.XI1.MM2 N_XI0.NET288_XI0.XI167.XI0.XI1.MM2_d
+ N_XI0.XI167.XI0.NET12_XI0.XI167.XI0.XI1.MM2_g N_VSS_XI0.XI167.XI0.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI0.XI166.XI0.XI1.MM2 N_XI0.NET282_XI0.XI166.XI0.XI1.MM2_d
+ N_XI0.XI166.XI0.NET12_XI0.XI166.XI0.XI1.MM2_g N_VSS_XI0.XI166.XI0.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI0.XI165.XI0.XI1.MM2 N_XI0.NET276_XI0.XI165.XI0.XI1.MM2_d
+ N_XI0.XI165.XI0.NET12_XI0.XI165.XI0.XI1.MM2_g N_VSS_XI0.XI165.XI0.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI0.XI159.XI0.XI1.MM2 N_XI0.NET270_XI0.XI159.XI0.XI1.MM2_d
+ N_XI0.XI159.XI0.NET12_XI0.XI159.XI0.XI1.MM2_g N_VSS_XI0.XI159.XI0.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI0.XI160.XI0.XI1.MM2 N_XI0.NET246_XI0.XI160.XI0.XI1.MM2_d
+ N_XI0.XI160.XI0.NET12_XI0.XI160.XI0.XI1.MM2_g N_VSS_XI0.XI160.XI0.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI0.XI161.XI0.XI1.MM2 N_XI0.NET252_XI0.XI161.XI0.XI1.MM2_d
+ N_XI0.XI161.XI0.NET12_XI0.XI161.XI0.XI1.MM2_g N_VSS_XI0.XI161.XI0.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI0.XI162.XI0.XI1.MM2 N_XI0.NET258_XI0.XI162.XI0.XI1.MM2_d
+ N_XI0.XI162.XI0.NET12_XI0.XI162.XI0.XI1.MM2_g N_VSS_XI0.XI162.XI0.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI0.XI121.XI0.XI1.MM2 N_XI0.NET264_XI0.XI121.XI0.XI1.MM2_d
+ N_XI0.XI121.XI0.NET12_XI0.XI121.XI0.XI1.MM2_g N_VSS_XI0.XI121.XI0.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI0.XI120.XI0.XI1.MM2 N_XI0.NET204_XI0.XI120.XI0.XI1.MM2_d
+ N_XI0.XI120.XI0.NET12_XI0.XI120.XI0.XI1.MM2_g N_VSS_XI0.XI120.XI0.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI0.XI119.XI0.XI1.MM2 N_XI0.NET210_XI0.XI119.XI0.XI1.MM2_d
+ N_XI0.XI119.XI0.NET12_XI0.XI119.XI0.XI1.MM2_g N_VSS_XI0.XI119.XI0.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI0.XI118.XI0.XI1.MM2 N_XI0.NET216_XI0.XI118.XI0.XI1.MM2_d
+ N_XI0.XI118.XI0.NET12_XI0.XI118.XI0.XI1.MM2_g N_VSS_XI0.XI118.XI0.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI0.XI91.XI0.XI1.MM2 N_XI0.NET222_XI0.XI91.XI0.XI1.MM2_d
+ N_XI0.XI91.XI0.NET12_XI0.XI91.XI0.XI1.MM2_g N_VSS_XI0.XI91.XI0.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI0.XI90.XI0.XI1.MM2 N_XI0.NET228_XI0.XI90.XI0.XI1.MM2_d
+ N_XI0.XI90.XI0.NET12_XI0.XI90.XI0.XI1.MM2_g N_VSS_XI0.XI90.XI0.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI0.XI89.XI0.XI1.MM2 N_XI0.NET240_XI0.XI89.XI0.XI1.MM2_d
+ N_XI0.XI89.XI0.NET12_XI0.XI89.XI0.XI1.MM2_g N_VSS_XI0.XI89.XI0.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI18.XI18.MM2 N_NET241_XI18.XI18.MM2_d N_XI18.XI18.NET7_XI18.XI18.MM2_g
+ N_NET508_XI18.XI18.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=3.075e-13 PD=1.48e-06 PS=1.23e-06
mXI18.XI19.MM2 N_NET242_XI18.XI19.MM2_d N_XI18.XI19.NET7_XI18.XI19.MM2_g
+ N_NET509_XI18.XI19.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=3.075e-13 PD=1.48e-06 PS=1.23e-06
mXI18.XI17.MM2 N_NET243_XI18.XI17.MM2_d N_XI18.XI17.NET7_XI18.XI17.MM2_g
+ N_NET510_XI18.XI17.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=3.075e-13 PD=1.48e-06 PS=1.23e-06
mXI18.XI16.MM2 N_NET244_XI18.XI16.MM2_d N_XI18.XI16.NET7_XI18.XI16.MM2_g
+ N_NET511_XI18.XI16.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=3.075e-13 PD=1.48e-06 PS=1.23e-06
mXI18.XI21.MM2 N_NET245_XI18.XI21.MM2_d N_XI18.XI21.NET7_XI18.XI21.MM2_g
+ N_NET512_XI18.XI21.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=3.075e-13 PD=1.48e-06 PS=1.23e-06
mXI18.XI20.MM2 N_NET246_XI18.XI20.MM2_d N_XI18.XI20.NET7_XI18.XI20.MM2_g
+ N_NET513_XI18.XI20.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=3.075e-13 PD=1.48e-06 PS=1.23e-06
mXI18.XI22.MM2 N_NET247_XI18.XI22.MM2_d N_XI18.XI22.NET7_XI18.XI22.MM2_g
+ N_NET514_XI18.XI22.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=3.075e-13 PD=1.48e-06 PS=1.23e-06
mXI18.XI6.MM2 N_NET248_XI18.XI6.MM2_d N_XI18.XI6.NET7_XI18.XI6.MM2_g
+ N_NET515_XI18.XI6.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=3.075e-13 PD=1.48e-06 PS=1.23e-06
mXI18.XI5.MM2 N_NET249_XI18.XI5.MM2_d N_XI18.XI5.NET7_XI18.XI5.MM2_g
+ N_NET516_XI18.XI5.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=3.075e-13 PD=1.48e-06 PS=1.23e-06
mXI18.XI7.MM2 N_NET250_XI18.XI7.MM2_d N_XI18.XI7.NET7_XI18.XI7.MM2_g
+ N_NET517_XI18.XI7.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=3.075e-13 PD=1.48e-06 PS=1.23e-06
mXI18.XI8.MM2 N_NET251_XI18.XI8.MM2_d N_XI18.XI8.NET7_XI18.XI8.MM2_g
+ N_NET518_XI18.XI8.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=3.075e-13 PD=1.48e-06 PS=1.23e-06
mXI18.XI3.MM2 N_NET252_XI18.XI3.MM2_d N_XI18.XI3.NET7_XI18.XI3.MM2_g
+ N_NET519_XI18.XI3.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=3.075e-13 PD=1.48e-06 PS=1.23e-06
mXI18.XI4.MM2 N_NET253_XI18.XI4.MM2_d N_XI18.XI4.NET7_XI18.XI4.MM2_g
+ N_NET520_XI18.XI4.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=3.075e-13 PD=1.48e-06 PS=1.23e-06
mXI18.XI2.MM2 N_NET254_XI18.XI2.MM2_d N_XI18.XI2.NET7_XI18.XI2.MM2_g
+ N_NET521_XI18.XI2.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=3.075e-13 PD=1.48e-06 PS=1.23e-06
mXI18.XI1.MM2 N_NET255_XI18.XI1.MM2_d N_XI18.XI1.NET7_XI18.XI1.MM2_g
+ N_NET522_XI18.XI1.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=3.075e-13 PD=1.48e-06 PS=1.23e-06
mXI18.XI0.MM2 N_NET256_XI18.XI0.MM2_d N_XI18.XI0.NET7_XI18.XI0.MM2_g
+ N_NET523_XI18.XI0.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=3.075e-13 PD=1.48e-06 PS=1.23e-06
mXI18.XI18.MM3 N_MIN15_XI18.XI18.MM3_d N_NET0859_XI18.XI18.MM3_g
+ N_NET508_XI18.XI18.MM3_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=6.05e-13 AS=3.075e-13 PD=2.92e-06 PS=1.23e-06
mXI18.XI19.MM3 N_MIN14_XI18.XI19.MM3_d N_NET0859_XI18.XI19.MM3_g
+ N_NET509_XI18.XI19.MM3_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=6.05e-13 AS=3.075e-13 PD=2.92e-06 PS=1.23e-06
mXI18.XI17.MM3 N_MIN13_XI18.XI17.MM3_d N_NET0859_XI18.XI17.MM3_g
+ N_NET510_XI18.XI17.MM3_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=6.05e-13 AS=3.075e-13 PD=2.92e-06 PS=1.23e-06
mXI18.XI16.MM3 N_MIN12_XI18.XI16.MM3_d N_NET0859_XI18.XI16.MM3_g
+ N_NET511_XI18.XI16.MM3_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=6.05e-13 AS=3.075e-13 PD=2.92e-06 PS=1.23e-06
mXI18.XI21.MM3 N_MIN11_XI18.XI21.MM3_d N_NET0859_XI18.XI21.MM3_g
+ N_NET512_XI18.XI21.MM3_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=6.05e-13 AS=3.075e-13 PD=2.92e-06 PS=1.23e-06
mXI18.XI20.MM3 N_MIN10_XI18.XI20.MM3_d N_NET0859_XI18.XI20.MM3_g
+ N_NET513_XI18.XI20.MM3_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=6.05e-13 AS=3.075e-13 PD=2.92e-06 PS=1.23e-06
mXI18.XI22.MM3 N_MIN9_XI18.XI22.MM3_d N_NET0859_XI18.XI22.MM3_g
+ N_NET514_XI18.XI22.MM3_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=6.05e-13 AS=3.075e-13 PD=2.92e-06 PS=1.23e-06
mXI18.XI6.MM3 N_MIN8_XI18.XI6.MM3_d N_NET0859_XI18.XI6.MM3_g
+ N_NET515_XI18.XI6.MM3_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=6.05e-13 AS=3.075e-13 PD=2.92e-06 PS=1.23e-06
mXI18.XI5.MM3 N_MIN7_XI18.XI5.MM3_d N_NET0859_XI18.XI5.MM3_g
+ N_NET516_XI18.XI5.MM3_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=6.05e-13 AS=3.075e-13 PD=2.92e-06 PS=1.23e-06
mXI18.XI7.MM3 N_MIN6_XI18.XI7.MM3_d N_NET0859_XI18.XI7.MM3_g
+ N_NET517_XI18.XI7.MM3_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=6.05e-13 AS=3.075e-13 PD=2.92e-06 PS=1.23e-06
mXI18.XI8.MM3 N_MIN5_XI18.XI8.MM3_d N_NET0859_XI18.XI8.MM3_g
+ N_NET518_XI18.XI8.MM3_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=6.05e-13 AS=3.075e-13 PD=2.92e-06 PS=1.23e-06
mXI18.XI3.MM3 N_MIN4_XI18.XI3.MM3_d N_NET0859_XI18.XI3.MM3_g
+ N_NET519_XI18.XI3.MM3_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=6.05e-13 AS=3.075e-13 PD=2.92e-06 PS=1.23e-06
mXI18.XI4.MM3 N_MIN3_XI18.XI4.MM3_d N_NET0859_XI18.XI4.MM3_g
+ N_NET520_XI18.XI4.MM3_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=6.05e-13 AS=3.075e-13 PD=2.92e-06 PS=1.23e-06
mXI18.XI2.MM3 N_MIN2_XI18.XI2.MM3_d N_NET0859_XI18.XI2.MM3_g
+ N_NET521_XI18.XI2.MM3_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=6.05e-13 AS=3.075e-13 PD=2.92e-06 PS=1.23e-06
mXI18.XI1.MM3 N_MIN1_XI18.XI1.MM3_d N_NET0859_XI18.XI1.MM3_g
+ N_NET522_XI18.XI1.MM3_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=6.05e-13 AS=3.075e-13 PD=2.92e-06 PS=1.23e-06
mXI18.XI0.MM3 N_MIN0_XI18.XI0.MM3_d N_NET0859_XI18.XI0.MM3_g
+ N_NET523_XI18.XI0.MM3_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=6.05e-13 AS=3.075e-13 PD=2.92e-06 PS=1.23e-06
mXI18.XI18.MM4 N_XI18.XI18.NET7_XI18.XI18.MM4_d N_NET0859_XI18.XI18.MM4_g
+ N_VSS_XI18.XI18.MM4_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI18.XI19.MM4 N_XI18.XI19.NET7_XI18.XI19.MM4_d N_NET0859_XI18.XI19.MM4_g
+ N_VSS_XI18.XI19.MM4_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI18.XI17.MM4 N_XI18.XI17.NET7_XI18.XI17.MM4_d N_NET0859_XI18.XI17.MM4_g
+ N_VSS_XI18.XI17.MM4_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI18.XI16.MM4 N_XI18.XI16.NET7_XI18.XI16.MM4_d N_NET0859_XI18.XI16.MM4_g
+ N_VSS_XI18.XI16.MM4_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI18.XI21.MM4 N_XI18.XI21.NET7_XI18.XI21.MM4_d N_NET0859_XI18.XI21.MM4_g
+ N_VSS_XI18.XI21.MM4_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI18.XI20.MM4 N_XI18.XI20.NET7_XI18.XI20.MM4_d N_NET0859_XI18.XI20.MM4_g
+ N_VSS_XI18.XI20.MM4_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI18.XI22.MM4 N_XI18.XI22.NET7_XI18.XI22.MM4_d N_NET0859_XI18.XI22.MM4_g
+ N_VSS_XI18.XI22.MM4_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI18.XI6.MM4 N_XI18.XI6.NET7_XI18.XI6.MM4_d N_NET0859_XI18.XI6.MM4_g
+ N_VSS_XI18.XI6.MM4_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI18.XI5.MM4 N_XI18.XI5.NET7_XI18.XI5.MM4_d N_NET0859_XI18.XI5.MM4_g
+ N_VSS_XI18.XI5.MM4_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI18.XI7.MM4 N_XI18.XI7.NET7_XI18.XI7.MM4_d N_NET0859_XI18.XI7.MM4_g
+ N_VSS_XI18.XI7.MM4_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI18.XI8.MM4 N_XI18.XI8.NET7_XI18.XI8.MM4_d N_NET0859_XI18.XI8.MM4_g
+ N_VSS_XI18.XI8.MM4_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI18.XI3.MM4 N_XI18.XI3.NET7_XI18.XI3.MM4_d N_NET0859_XI18.XI3.MM4_g
+ N_VSS_XI18.XI3.MM4_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI18.XI4.MM4 N_XI18.XI4.NET7_XI18.XI4.MM4_d N_NET0859_XI18.XI4.MM4_g
+ N_VSS_XI18.XI4.MM4_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI18.XI2.MM4 N_XI18.XI2.NET7_XI18.XI2.MM4_d N_NET0859_XI18.XI2.MM4_g
+ N_VSS_XI18.XI2.MM4_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI18.XI1.MM4 N_XI18.XI1.NET7_XI18.XI1.MM4_d N_NET0859_XI18.XI1.MM4_g
+ N_VSS_XI18.XI1.MM4_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI18.XI0.MM4 N_XI18.XI0.NET7_XI18.XI0.MM4_d N_NET0859_XI18.XI0.MM4_g
+ N_VSS_XI18.XI0.MM4_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI15.MM1 N_XI15.NET40_XI15.MM1_d N_NET198_XI15.MM1_g N_VSS_XI15.MM1_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI15.XI16.XI1.MM2 N_XI15.XI16.XI1.NET036_XI15.XI16.XI1.MM2_d
+ N_NET198_XI15.XI16.XI1.MM2_g N_VSS_XI15.XI16.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.375e-13 AS=2.45e-13
+ PD=5.5e-07 PS=1.48e-06
mXI15.XI16.XI1.MM0 N_XI15.XI16.NET6_XI15.XI16.XI1.MM0_d
+ N_NET508_XI15.XI16.XI1.MM0_g N_XI15.XI16.XI1.NET036_XI15.XI16.XI1.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=1.375e-13
+ PD=1.52e-06 PS=5.5e-07
mXI15.XI16.XI0.MM2 N_NET417_XI15.XI16.XI0.MM2_d
+ N_XI15.XI16.NET6_XI15.XI16.XI0.MM2_g N_VSS_XI15.XI16.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI15.XI17.XI0.MM2 N_XI15.XI17.NET12_XI15.XI17.XI0.MM2_d
+ N_XI15.NET40_XI15.XI17.XI0.MM2_g N_VSS_XI15.XI17.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.875e-13 AS=2.45e-13
+ PD=7.5e-07 PS=1.48e-06
mXI15.XI17.XI0.MM0 N_XI15.XI17.NET12_XI15.XI17.XI0.MM0_d
+ N_NET509_XI15.XI17.XI0.MM0_g N_VSS_XI15.XI17.XI0.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.875e-13 AS=2.55e-13
+ PD=7.5e-07 PS=1.52e-06
mXI15.XI17.XI1.MM2 N_NET418_XI15.XI17.XI1.MM2_d
+ N_XI15.XI17.NET12_XI15.XI17.XI1.MM2_g N_VSS_XI15.XI17.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI15.XI18.XI0.MM2 N_XI15.XI18.NET12_XI15.XI18.XI0.MM2_d
+ N_XI15.NET40_XI15.XI18.XI0.MM2_g N_VSS_XI15.XI18.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.875e-13 AS=2.45e-13
+ PD=7.5e-07 PS=1.48e-06
mXI15.XI18.XI0.MM0 N_XI15.XI18.NET12_XI15.XI18.XI0.MM0_d
+ N_NET510_XI15.XI18.XI0.MM0_g N_VSS_XI15.XI18.XI0.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.875e-13 AS=2.55e-13
+ PD=7.5e-07 PS=1.52e-06
mXI15.XI18.XI1.MM2 N_NET419_XI15.XI18.XI1.MM2_d
+ N_XI15.XI18.NET12_XI15.XI18.XI1.MM2_g N_VSS_XI15.XI18.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI15.XI19.XI0.MM2 N_XI15.XI19.NET12_XI15.XI19.XI0.MM2_d
+ N_XI15.NET40_XI15.XI19.XI0.MM2_g N_VSS_XI15.XI19.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.875e-13 AS=2.45e-13
+ PD=7.5e-07 PS=1.48e-06
mXI15.XI19.XI0.MM0 N_XI15.XI19.NET12_XI15.XI19.XI0.MM0_d
+ N_NET511_XI15.XI19.XI0.MM0_g N_VSS_XI15.XI19.XI0.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.875e-13 AS=2.55e-13
+ PD=7.5e-07 PS=1.52e-06
mXI15.XI19.XI1.MM2 N_NET420_XI15.XI19.XI1.MM2_d
+ N_XI15.XI19.NET12_XI15.XI19.XI1.MM2_g N_VSS_XI15.XI19.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI15.XI20.XI0.MM2 N_XI15.XI20.NET12_XI15.XI20.XI0.MM2_d
+ N_XI15.NET40_XI15.XI20.XI0.MM2_g N_VSS_XI15.XI20.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.875e-13 AS=2.45e-13
+ PD=7.5e-07 PS=1.48e-06
mXI15.XI20.XI0.MM0 N_XI15.XI20.NET12_XI15.XI20.XI0.MM0_d
+ N_NET512_XI15.XI20.XI0.MM0_g N_VSS_XI15.XI20.XI0.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.875e-13 AS=2.55e-13
+ PD=7.5e-07 PS=1.52e-06
mXI15.XI20.XI1.MM2 N_NET421_XI15.XI20.XI1.MM2_d
+ N_XI15.XI20.NET12_XI15.XI20.XI1.MM2_g N_VSS_XI15.XI20.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI15.XI21.XI0.MM2 N_XI15.XI21.NET12_XI15.XI21.XI0.MM2_d
+ N_XI15.NET40_XI15.XI21.XI0.MM2_g N_VSS_XI15.XI21.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.875e-13 AS=2.45e-13
+ PD=7.5e-07 PS=1.48e-06
mXI15.XI21.XI0.MM0 N_XI15.XI21.NET12_XI15.XI21.XI0.MM0_d
+ N_NET513_XI15.XI21.XI0.MM0_g N_VSS_XI15.XI21.XI0.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.875e-13 AS=2.55e-13
+ PD=7.5e-07 PS=1.52e-06
mXI15.XI21.XI1.MM2 N_NET422_XI15.XI21.XI1.MM2_d
+ N_XI15.XI21.NET12_XI15.XI21.XI1.MM2_g N_VSS_XI15.XI21.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI15.XI22.XI0.MM2 N_XI15.XI22.NET12_XI15.XI22.XI0.MM2_d
+ N_XI15.NET40_XI15.XI22.XI0.MM2_g N_VSS_XI15.XI22.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.875e-13 AS=2.45e-13
+ PD=7.5e-07 PS=1.48e-06
mXI15.XI22.XI0.MM0 N_XI15.XI22.NET12_XI15.XI22.XI0.MM0_d
+ N_NET514_XI15.XI22.XI0.MM0_g N_VSS_XI15.XI22.XI0.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.875e-13 AS=2.55e-13
+ PD=7.5e-07 PS=1.52e-06
mXI15.XI22.XI1.MM2 N_NET423_XI15.XI22.XI1.MM2_d
+ N_XI15.XI22.NET12_XI15.XI22.XI1.MM2_g N_VSS_XI15.XI22.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI15.XI23.XI0.MM2 N_XI15.XI23.NET12_XI15.XI23.XI0.MM2_d
+ N_XI15.NET40_XI15.XI23.XI0.MM2_g N_VSS_XI15.XI23.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.875e-13 AS=2.45e-13
+ PD=7.5e-07 PS=1.48e-06
mXI15.XI23.XI0.MM0 N_XI15.XI23.NET12_XI15.XI23.XI0.MM0_d
+ N_NET515_XI15.XI23.XI0.MM0_g N_VSS_XI15.XI23.XI0.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.875e-13 AS=2.55e-13
+ PD=7.5e-07 PS=1.52e-06
mXI15.XI23.XI1.MM2 N_NET424_XI15.XI23.XI1.MM2_d
+ N_XI15.XI23.NET12_XI15.XI23.XI1.MM2_g N_VSS_XI15.XI23.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI15.XI24.XI0.MM2 N_XI15.XI24.NET12_XI15.XI24.XI0.MM2_d
+ N_XI15.NET40_XI15.XI24.XI0.MM2_g N_VSS_XI15.XI24.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.875e-13 AS=2.45e-13
+ PD=7.5e-07 PS=1.48e-06
mXI15.XI24.XI0.MM0 N_XI15.XI24.NET12_XI15.XI24.XI0.MM0_d
+ N_NET516_XI15.XI24.XI0.MM0_g N_VSS_XI15.XI24.XI0.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.875e-13 AS=2.55e-13
+ PD=7.5e-07 PS=1.52e-06
mXI15.XI24.XI1.MM2 N_NET425_XI15.XI24.XI1.MM2_d
+ N_XI15.XI24.NET12_XI15.XI24.XI1.MM2_g N_VSS_XI15.XI24.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI15.XI25.XI0.MM2 N_XI15.XI25.NET12_XI15.XI25.XI0.MM2_d
+ N_XI15.NET40_XI15.XI25.XI0.MM2_g N_VSS_XI15.XI25.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.875e-13 AS=2.45e-13
+ PD=7.5e-07 PS=1.48e-06
mXI15.XI25.XI0.MM0 N_XI15.XI25.NET12_XI15.XI25.XI0.MM0_d
+ N_NET517_XI15.XI25.XI0.MM0_g N_VSS_XI15.XI25.XI0.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.875e-13 AS=2.55e-13
+ PD=7.5e-07 PS=1.52e-06
mXI15.XI25.XI1.MM2 N_NET426_XI15.XI25.XI1.MM2_d
+ N_XI15.XI25.NET12_XI15.XI25.XI1.MM2_g N_VSS_XI15.XI25.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI15.XI26.XI0.MM2 N_XI15.XI26.NET12_XI15.XI26.XI0.MM2_d
+ N_XI15.NET40_XI15.XI26.XI0.MM2_g N_VSS_XI15.XI26.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.875e-13 AS=2.45e-13
+ PD=7.5e-07 PS=1.48e-06
mXI15.XI26.XI0.MM0 N_XI15.XI26.NET12_XI15.XI26.XI0.MM0_d
+ N_NET518_XI15.XI26.XI0.MM0_g N_VSS_XI15.XI26.XI0.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.875e-13 AS=2.55e-13
+ PD=7.5e-07 PS=1.52e-06
mXI15.XI26.XI1.MM2 N_NET427_XI15.XI26.XI1.MM2_d
+ N_XI15.XI26.NET12_XI15.XI26.XI1.MM2_g N_VSS_XI15.XI26.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI15.XI27.XI0.MM2 N_XI15.XI27.NET12_XI15.XI27.XI0.MM2_d
+ N_XI15.NET40_XI15.XI27.XI0.MM2_g N_VSS_XI15.XI27.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.875e-13 AS=2.45e-13
+ PD=7.5e-07 PS=1.48e-06
mXI15.XI27.XI0.MM0 N_XI15.XI27.NET12_XI15.XI27.XI0.MM0_d
+ N_NET519_XI15.XI27.XI0.MM0_g N_VSS_XI15.XI27.XI0.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.875e-13 AS=2.55e-13
+ PD=7.5e-07 PS=1.52e-06
mXI15.XI27.XI1.MM2 N_NET428_XI15.XI27.XI1.MM2_d
+ N_XI15.XI27.NET12_XI15.XI27.XI1.MM2_g N_VSS_XI15.XI27.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI15.XI28.XI0.MM2 N_XI15.XI28.NET12_XI15.XI28.XI0.MM2_d
+ N_XI15.NET40_XI15.XI28.XI0.MM2_g N_VSS_XI15.XI28.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.875e-13 AS=2.45e-13
+ PD=7.5e-07 PS=1.48e-06
mXI15.XI28.XI0.MM0 N_XI15.XI28.NET12_XI15.XI28.XI0.MM0_d
+ N_NET520_XI15.XI28.XI0.MM0_g N_VSS_XI15.XI28.XI0.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.875e-13 AS=2.55e-13
+ PD=7.5e-07 PS=1.52e-06
mXI15.XI28.XI1.MM2 N_NET429_XI15.XI28.XI1.MM2_d
+ N_XI15.XI28.NET12_XI15.XI28.XI1.MM2_g N_VSS_XI15.XI28.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI15.XI29.XI0.MM2 N_XI15.XI29.NET12_XI15.XI29.XI0.MM2_d
+ N_XI15.NET40_XI15.XI29.XI0.MM2_g N_VSS_XI15.XI29.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.875e-13 AS=2.45e-13
+ PD=7.5e-07 PS=1.48e-06
mXI15.XI29.XI0.MM0 N_XI15.XI29.NET12_XI15.XI29.XI0.MM0_d
+ N_NET521_XI15.XI29.XI0.MM0_g N_VSS_XI15.XI29.XI0.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.875e-13 AS=2.55e-13
+ PD=7.5e-07 PS=1.52e-06
mXI15.XI29.XI1.MM2 N_NET430_XI15.XI29.XI1.MM2_d
+ N_XI15.XI29.NET12_XI15.XI29.XI1.MM2_g N_VSS_XI15.XI29.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI15.XI30.XI0.MM2 N_XI15.XI30.NET12_XI15.XI30.XI0.MM2_d
+ N_XI15.NET40_XI15.XI30.XI0.MM2_g N_VSS_XI15.XI30.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.875e-13 AS=2.45e-13
+ PD=7.5e-07 PS=1.48e-06
mXI15.XI30.XI0.MM0 N_XI15.XI30.NET12_XI15.XI30.XI0.MM0_d
+ N_NET522_XI15.XI30.XI0.MM0_g N_VSS_XI15.XI30.XI0.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.875e-13 AS=2.55e-13
+ PD=7.5e-07 PS=1.52e-06
mXI15.XI30.XI1.MM2 N_NET431_XI15.XI30.XI1.MM2_d
+ N_XI15.XI30.NET12_XI15.XI30.XI1.MM2_g N_VSS_XI15.XI30.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI15.XI31.XI0.MM2 N_XI15.XI31.NET12_XI15.XI31.XI0.MM2_d
+ N_XI15.NET40_XI15.XI31.XI0.MM2_g N_VSS_XI15.XI31.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.875e-13 AS=2.45e-13
+ PD=7.5e-07 PS=1.48e-06
mXI15.XI31.XI0.MM0 N_XI15.XI31.NET12_XI15.XI31.XI0.MM0_d
+ N_NET523_XI15.XI31.XI0.MM0_g N_VSS_XI15.XI31.XI0.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.875e-13 AS=2.55e-13
+ PD=7.5e-07 PS=1.52e-06
mXI15.XI31.XI1.MM2 N_NET432_XI15.XI31.XI1.MM2_d
+ N_XI15.XI31.NET12_XI15.XI31.XI1.MM2_g N_VSS_XI15.XI31.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI12.XI30.XI0.MM2 N_XI12.XI30.NET0180_XI12.XI30.XI0.MM2_d
+ N_NET222_XI12.XI30.XI0.MM2_g N_VSS_XI12.XI30.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI29.XI0.MM2 N_XI12.XI29.NET0180_XI12.XI29.XI0.MM2_d
+ N_NET222_XI12.XI29.XI0.MM2_g N_VSS_XI12.XI29.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI31.XI0.MM2 N_XI12.XI31.NET0180_XI12.XI31.XI0.MM2_d
+ N_NET222_XI12.XI31.XI0.MM2_g N_VSS_XI12.XI31.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI28.XI0.MM2 N_XI12.XI28.NET0180_XI12.XI28.XI0.MM2_d
+ N_NET222_XI12.XI28.XI0.MM2_g N_VSS_XI12.XI28.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI25.XI0.MM2 N_XI12.XI25.NET0180_XI12.XI25.XI0.MM2_d
+ N_NET222_XI12.XI25.XI0.MM2_g N_VSS_XI12.XI25.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI26.XI0.MM2 N_XI12.XI26.NET0180_XI12.XI26.XI0.MM2_d
+ N_NET222_XI12.XI26.XI0.MM2_g N_VSS_XI12.XI26.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI24.XI0.MM2 N_XI12.XI24.NET0180_XI12.XI24.XI0.MM2_d
+ N_NET222_XI12.XI24.XI0.MM2_g N_VSS_XI12.XI24.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI27.XI0.MM2 N_XI12.XI27.NET0180_XI12.XI27.XI0.MM2_d
+ N_NET222_XI12.XI27.XI0.MM2_g N_VSS_XI12.XI27.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI22.XI0.MM2 N_XI12.XI22.NET0180_XI12.XI22.XI0.MM2_d
+ N_NET222_XI12.XI22.XI0.MM2_g N_VSS_XI12.XI22.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI21.XI0.MM2 N_XI12.XI21.NET0180_XI12.XI21.XI0.MM2_d
+ N_NET222_XI12.XI21.XI0.MM2_g N_VSS_XI12.XI21.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI23.XI0.MM2 N_XI12.XI23.NET0180_XI12.XI23.XI0.MM2_d
+ N_NET222_XI12.XI23.XI0.MM2_g N_VSS_XI12.XI23.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI19.XI0.MM2 N_XI12.XI19.NET0180_XI12.XI19.XI0.MM2_d
+ N_NET222_XI12.XI19.XI0.MM2_g N_VSS_XI12.XI19.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI20.XI0.MM2 N_XI12.XI20.NET0180_XI12.XI20.XI0.MM2_d
+ N_NET222_XI12.XI20.XI0.MM2_g N_VSS_XI12.XI20.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI18.XI0.MM2 N_XI12.XI18.NET0180_XI12.XI18.XI0.MM2_d
+ N_NET222_XI12.XI18.XI0.MM2_g N_VSS_XI12.XI18.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI17.XI0.MM2 N_XI12.XI17.NET0180_XI12.XI17.XI0.MM2_d
+ N_NET222_XI12.XI17.XI0.MM2_g N_VSS_XI12.XI17.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI0.XI0.MM2 N_XI12.XI0.NET0180_XI12.XI0.XI0.MM2_d
+ N_NET222_XI12.XI0.XI0.MM2_g N_VSS_XI12.XI0.XI0.MM2_s N_VSS_XI10.XI0.XI0.MM2_b
+ N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI12.XI30.XI1.MM2 N_XI12.XI30.NET35_XI12.XI30.XI1.MM2_d
+ N_XI12.XI30.NET0180_XI12.XI30.XI1.MM2_g N_VSS_XI12.XI30.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI29.XI1.MM2 N_XI12.XI29.NET35_XI12.XI29.XI1.MM2_d
+ N_XI12.XI29.NET0180_XI12.XI29.XI1.MM2_g N_VSS_XI12.XI29.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI31.XI1.MM2 N_XI12.XI31.NET35_XI12.XI31.XI1.MM2_d
+ N_XI12.XI31.NET0180_XI12.XI31.XI1.MM2_g N_VSS_XI12.XI31.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI28.XI1.MM2 N_XI12.XI28.NET35_XI12.XI28.XI1.MM2_d
+ N_XI12.XI28.NET0180_XI12.XI28.XI1.MM2_g N_VSS_XI12.XI28.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI25.XI1.MM2 N_XI12.XI25.NET35_XI12.XI25.XI1.MM2_d
+ N_XI12.XI25.NET0180_XI12.XI25.XI1.MM2_g N_VSS_XI12.XI25.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI26.XI1.MM2 N_XI12.XI26.NET35_XI12.XI26.XI1.MM2_d
+ N_XI12.XI26.NET0180_XI12.XI26.XI1.MM2_g N_VSS_XI12.XI26.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI24.XI1.MM2 N_XI12.XI24.NET35_XI12.XI24.XI1.MM2_d
+ N_XI12.XI24.NET0180_XI12.XI24.XI1.MM2_g N_VSS_XI12.XI24.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI27.XI1.MM2 N_XI12.XI27.NET35_XI12.XI27.XI1.MM2_d
+ N_XI12.XI27.NET0180_XI12.XI27.XI1.MM2_g N_VSS_XI12.XI27.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI22.XI1.MM2 N_XI12.XI22.NET35_XI12.XI22.XI1.MM2_d
+ N_XI12.XI22.NET0180_XI12.XI22.XI1.MM2_g N_VSS_XI12.XI22.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI21.XI1.MM2 N_XI12.XI21.NET35_XI12.XI21.XI1.MM2_d
+ N_XI12.XI21.NET0180_XI12.XI21.XI1.MM2_g N_VSS_XI12.XI21.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI23.XI1.MM2 N_XI12.XI23.NET35_XI12.XI23.XI1.MM2_d
+ N_XI12.XI23.NET0180_XI12.XI23.XI1.MM2_g N_VSS_XI12.XI23.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI19.XI1.MM2 N_XI12.XI19.NET35_XI12.XI19.XI1.MM2_d
+ N_XI12.XI19.NET0180_XI12.XI19.XI1.MM2_g N_VSS_XI12.XI19.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI20.XI1.MM2 N_XI12.XI20.NET35_XI12.XI20.XI1.MM2_d
+ N_XI12.XI20.NET0180_XI12.XI20.XI1.MM2_g N_VSS_XI12.XI20.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI18.XI1.MM2 N_XI12.XI18.NET35_XI12.XI18.XI1.MM2_d
+ N_XI12.XI18.NET0180_XI12.XI18.XI1.MM2_g N_VSS_XI12.XI18.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI17.XI1.MM2 N_XI12.XI17.NET35_XI12.XI17.XI1.MM2_d
+ N_XI12.XI17.NET0180_XI12.XI17.XI1.MM2_g N_VSS_XI12.XI17.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI0.XI1.MM2 N_XI12.XI0.NET35_XI12.XI0.XI1.MM2_d
+ N_XI12.XI0.NET0180_XI12.XI0.XI1.MM2_g N_VSS_XI12.XI0.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI30.MM26 N_XI12.XI30.CLKB_XI12.XI30.MM26_d
+ N_XI12.XI30.NET35_XI12.XI30.MM26_g N_VSS_XI12.XI30.MM26_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI29.MM26 N_XI12.XI29.CLKB_XI12.XI29.MM26_d
+ N_XI12.XI29.NET35_XI12.XI29.MM26_g N_VSS_XI12.XI29.MM26_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI31.MM26 N_XI12.XI31.CLKB_XI12.XI31.MM26_d
+ N_XI12.XI31.NET35_XI12.XI31.MM26_g N_VSS_XI12.XI31.MM26_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI28.MM26 N_XI12.XI28.CLKB_XI12.XI28.MM26_d
+ N_XI12.XI28.NET35_XI12.XI28.MM26_g N_VSS_XI12.XI28.MM26_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI25.MM26 N_XI12.XI25.CLKB_XI12.XI25.MM26_d
+ N_XI12.XI25.NET35_XI12.XI25.MM26_g N_VSS_XI12.XI25.MM26_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI26.MM26 N_XI12.XI26.CLKB_XI12.XI26.MM26_d
+ N_XI12.XI26.NET35_XI12.XI26.MM26_g N_VSS_XI12.XI26.MM26_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI24.MM26 N_XI12.XI24.CLKB_XI12.XI24.MM26_d
+ N_XI12.XI24.NET35_XI12.XI24.MM26_g N_VSS_XI12.XI24.MM26_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI27.MM26 N_XI12.XI27.CLKB_XI12.XI27.MM26_d
+ N_XI12.XI27.NET35_XI12.XI27.MM26_g N_VSS_XI12.XI27.MM26_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI22.MM26 N_XI12.XI22.CLKB_XI12.XI22.MM26_d
+ N_XI12.XI22.NET35_XI12.XI22.MM26_g N_VSS_XI12.XI22.MM26_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI21.MM26 N_XI12.XI21.CLKB_XI12.XI21.MM26_d
+ N_XI12.XI21.NET35_XI12.XI21.MM26_g N_VSS_XI12.XI21.MM26_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI23.MM26 N_XI12.XI23.CLKB_XI12.XI23.MM26_d
+ N_XI12.XI23.NET35_XI12.XI23.MM26_g N_VSS_XI12.XI23.MM26_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI19.MM26 N_XI12.XI19.CLKB_XI12.XI19.MM26_d
+ N_XI12.XI19.NET35_XI12.XI19.MM26_g N_VSS_XI12.XI19.MM26_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI20.MM26 N_XI12.XI20.CLKB_XI12.XI20.MM26_d
+ N_XI12.XI20.NET35_XI12.XI20.MM26_g N_VSS_XI12.XI20.MM26_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI18.MM26 N_XI12.XI18.CLKB_XI12.XI18.MM26_d
+ N_XI12.XI18.NET35_XI12.XI18.MM26_g N_VSS_XI12.XI18.MM26_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI17.MM26 N_XI12.XI17.CLKB_XI12.XI17.MM26_d
+ N_XI12.XI17.NET35_XI12.XI17.MM26_g N_VSS_XI12.XI17.MM26_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI0.MM26 N_XI12.XI0.CLKB_XI12.XI0.MM26_d N_XI12.XI0.NET35_XI12.XI0.MM26_g
+ N_VSS_XI12.XI0.MM26_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI12.XI30.MM19 N_XI12.XI30.NET27_XI12.XI30.MM19_d N_NET417_XI12.XI30.MM19_g
+ N_VSS_XI12.XI30.MM19_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI12.XI29.MM19 N_XI12.XI29.NET27_XI12.XI29.MM19_d N_NET418_XI12.XI29.MM19_g
+ N_VSS_XI12.XI29.MM19_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI12.XI31.MM19 N_XI12.XI31.NET27_XI12.XI31.MM19_d N_NET419_XI12.XI31.MM19_g
+ N_VSS_XI12.XI31.MM19_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI12.XI28.MM19 N_XI12.XI28.NET27_XI12.XI28.MM19_d N_NET420_XI12.XI28.MM19_g
+ N_VSS_XI12.XI28.MM19_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI12.XI25.MM19 N_XI12.XI25.NET27_XI12.XI25.MM19_d N_NET421_XI12.XI25.MM19_g
+ N_VSS_XI12.XI25.MM19_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI12.XI26.MM19 N_XI12.XI26.NET27_XI12.XI26.MM19_d N_NET422_XI12.XI26.MM19_g
+ N_VSS_XI12.XI26.MM19_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI12.XI24.MM19 N_XI12.XI24.NET27_XI12.XI24.MM19_d N_NET423_XI12.XI24.MM19_g
+ N_VSS_XI12.XI24.MM19_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI12.XI27.MM19 N_XI12.XI27.NET27_XI12.XI27.MM19_d N_NET424_XI12.XI27.MM19_g
+ N_VSS_XI12.XI27.MM19_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI12.XI22.MM19 N_XI12.XI22.NET27_XI12.XI22.MM19_d N_NET425_XI12.XI22.MM19_g
+ N_VSS_XI12.XI22.MM19_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI12.XI21.MM19 N_XI12.XI21.NET27_XI12.XI21.MM19_d N_NET426_XI12.XI21.MM19_g
+ N_VSS_XI12.XI21.MM19_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI12.XI23.MM19 N_XI12.XI23.NET27_XI12.XI23.MM19_d N_NET427_XI12.XI23.MM19_g
+ N_VSS_XI12.XI23.MM19_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI12.XI19.MM19 N_XI12.XI19.NET27_XI12.XI19.MM19_d N_NET428_XI12.XI19.MM19_g
+ N_VSS_XI12.XI19.MM19_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI12.XI20.MM19 N_XI12.XI20.NET27_XI12.XI20.MM19_d N_NET429_XI12.XI20.MM19_g
+ N_VSS_XI12.XI20.MM19_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI12.XI18.MM19 N_XI12.XI18.NET27_XI12.XI18.MM19_d N_NET430_XI12.XI18.MM19_g
+ N_VSS_XI12.XI18.MM19_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI12.XI17.MM19 N_XI12.XI17.NET27_XI12.XI17.MM19_d N_NET431_XI12.XI17.MM19_g
+ N_VSS_XI12.XI17.MM19_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI12.XI0.MM19 N_XI12.XI0.NET27_XI12.XI0.MM19_d N_NET432_XI12.XI0.MM19_g
+ N_VSS_XI12.XI0.MM19_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI12.XI30.MM18 N_XI12.XI30.NET31_XI12.XI30.MM18_d
+ N_XI12.XI30.NET27_XI12.XI30.MM18_g N_VSS_XI12.XI30.MM18_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI29.MM18 N_XI12.XI29.NET31_XI12.XI29.MM18_d
+ N_XI12.XI29.NET27_XI12.XI29.MM18_g N_VSS_XI12.XI29.MM18_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI31.MM18 N_XI12.XI31.NET31_XI12.XI31.MM18_d
+ N_XI12.XI31.NET27_XI12.XI31.MM18_g N_VSS_XI12.XI31.MM18_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI28.MM18 N_XI12.XI28.NET31_XI12.XI28.MM18_d
+ N_XI12.XI28.NET27_XI12.XI28.MM18_g N_VSS_XI12.XI28.MM18_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI25.MM18 N_XI12.XI25.NET31_XI12.XI25.MM18_d
+ N_XI12.XI25.NET27_XI12.XI25.MM18_g N_VSS_XI12.XI25.MM18_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI26.MM18 N_XI12.XI26.NET31_XI12.XI26.MM18_d
+ N_XI12.XI26.NET27_XI12.XI26.MM18_g N_VSS_XI12.XI26.MM18_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI24.MM18 N_XI12.XI24.NET31_XI12.XI24.MM18_d
+ N_XI12.XI24.NET27_XI12.XI24.MM18_g N_VSS_XI12.XI24.MM18_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI27.MM18 N_XI12.XI27.NET31_XI12.XI27.MM18_d
+ N_XI12.XI27.NET27_XI12.XI27.MM18_g N_VSS_XI12.XI27.MM18_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI22.MM18 N_XI12.XI22.NET31_XI12.XI22.MM18_d
+ N_XI12.XI22.NET27_XI12.XI22.MM18_g N_VSS_XI12.XI22.MM18_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI21.MM18 N_XI12.XI21.NET31_XI12.XI21.MM18_d
+ N_XI12.XI21.NET27_XI12.XI21.MM18_g N_VSS_XI12.XI21.MM18_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI23.MM18 N_XI12.XI23.NET31_XI12.XI23.MM18_d
+ N_XI12.XI23.NET27_XI12.XI23.MM18_g N_VSS_XI12.XI23.MM18_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI19.MM18 N_XI12.XI19.NET31_XI12.XI19.MM18_d
+ N_XI12.XI19.NET27_XI12.XI19.MM18_g N_VSS_XI12.XI19.MM18_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI20.MM18 N_XI12.XI20.NET31_XI12.XI20.MM18_d
+ N_XI12.XI20.NET27_XI12.XI20.MM18_g N_VSS_XI12.XI20.MM18_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI18.MM18 N_XI12.XI18.NET31_XI12.XI18.MM18_d
+ N_XI12.XI18.NET27_XI12.XI18.MM18_g N_VSS_XI12.XI18.MM18_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI17.MM18 N_XI12.XI17.NET31_XI12.XI17.MM18_d
+ N_XI12.XI17.NET27_XI12.XI17.MM18_g N_VSS_XI12.XI17.MM18_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI0.MM18 N_XI12.XI0.NET31_XI12.XI0.MM18_d N_XI12.XI0.NET27_XI12.XI0.MM18_g
+ N_VSS_XI12.XI0.MM18_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI12.XI30.MM28 N_XI12.XI30.NET31_XI12.XI30.MM28_d
+ N_XI12.XI30.CLKB_XI12.XI30.MM28_g N_XI12.XI30.NET58_XI12.XI30.MM28_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI29.MM28 N_XI12.XI29.NET31_XI12.XI29.MM28_d
+ N_XI12.XI29.CLKB_XI12.XI29.MM28_g N_XI12.XI29.NET58_XI12.XI29.MM28_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI31.MM28 N_XI12.XI31.NET31_XI12.XI31.MM28_d
+ N_XI12.XI31.CLKB_XI12.XI31.MM28_g N_XI12.XI31.NET58_XI12.XI31.MM28_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI28.MM28 N_XI12.XI28.NET31_XI12.XI28.MM28_d
+ N_XI12.XI28.CLKB_XI12.XI28.MM28_g N_XI12.XI28.NET58_XI12.XI28.MM28_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI25.MM28 N_XI12.XI25.NET31_XI12.XI25.MM28_d
+ N_XI12.XI25.CLKB_XI12.XI25.MM28_g N_XI12.XI25.NET58_XI12.XI25.MM28_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI26.MM28 N_XI12.XI26.NET31_XI12.XI26.MM28_d
+ N_XI12.XI26.CLKB_XI12.XI26.MM28_g N_XI12.XI26.NET58_XI12.XI26.MM28_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI24.MM28 N_XI12.XI24.NET31_XI12.XI24.MM28_d
+ N_XI12.XI24.CLKB_XI12.XI24.MM28_g N_XI12.XI24.NET58_XI12.XI24.MM28_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI27.MM28 N_XI12.XI27.NET31_XI12.XI27.MM28_d
+ N_XI12.XI27.CLKB_XI12.XI27.MM28_g N_XI12.XI27.NET58_XI12.XI27.MM28_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI22.MM28 N_XI12.XI22.NET31_XI12.XI22.MM28_d
+ N_XI12.XI22.CLKB_XI12.XI22.MM28_g N_XI12.XI22.NET58_XI12.XI22.MM28_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI21.MM28 N_XI12.XI21.NET31_XI12.XI21.MM28_d
+ N_XI12.XI21.CLKB_XI12.XI21.MM28_g N_XI12.XI21.NET58_XI12.XI21.MM28_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI23.MM28 N_XI12.XI23.NET31_XI12.XI23.MM28_d
+ N_XI12.XI23.CLKB_XI12.XI23.MM28_g N_XI12.XI23.NET58_XI12.XI23.MM28_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI19.MM28 N_XI12.XI19.NET31_XI12.XI19.MM28_d
+ N_XI12.XI19.CLKB_XI12.XI19.MM28_g N_XI12.XI19.NET58_XI12.XI19.MM28_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI20.MM28 N_XI12.XI20.NET31_XI12.XI20.MM28_d
+ N_XI12.XI20.CLKB_XI12.XI20.MM28_g N_XI12.XI20.NET58_XI12.XI20.MM28_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI18.MM28 N_XI12.XI18.NET31_XI12.XI18.MM28_d
+ N_XI12.XI18.CLKB_XI12.XI18.MM28_g N_XI12.XI18.NET58_XI12.XI18.MM28_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI17.MM28 N_XI12.XI17.NET31_XI12.XI17.MM28_d
+ N_XI12.XI17.CLKB_XI12.XI17.MM28_g N_XI12.XI17.NET58_XI12.XI17.MM28_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI0.MM28 N_XI12.XI0.NET31_XI12.XI0.MM28_d N_XI12.XI0.CLKB_XI12.XI0.MM28_g
+ N_XI12.XI0.NET58_XI12.XI0.MM28_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI12.XI30.MM6 N_XI12.XI30.NET15_XI12.XI30.MM6_d
+ N_XI12.XI30.NET58_XI12.XI30.MM6_g N_VSS_XI12.XI30.MM6_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI29.MM6 N_XI12.XI29.NET15_XI12.XI29.MM6_d
+ N_XI12.XI29.NET58_XI12.XI29.MM6_g N_VSS_XI12.XI29.MM6_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI31.MM6 N_XI12.XI31.NET15_XI12.XI31.MM6_d
+ N_XI12.XI31.NET58_XI12.XI31.MM6_g N_VSS_XI12.XI31.MM6_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI28.MM6 N_XI12.XI28.NET15_XI12.XI28.MM6_d
+ N_XI12.XI28.NET58_XI12.XI28.MM6_g N_VSS_XI12.XI28.MM6_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI25.MM6 N_XI12.XI25.NET15_XI12.XI25.MM6_d
+ N_XI12.XI25.NET58_XI12.XI25.MM6_g N_VSS_XI12.XI25.MM6_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI26.MM6 N_XI12.XI26.NET15_XI12.XI26.MM6_d
+ N_XI12.XI26.NET58_XI12.XI26.MM6_g N_VSS_XI12.XI26.MM6_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI24.MM6 N_XI12.XI24.NET15_XI12.XI24.MM6_d
+ N_XI12.XI24.NET58_XI12.XI24.MM6_g N_VSS_XI12.XI24.MM6_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI27.MM6 N_XI12.XI27.NET15_XI12.XI27.MM6_d
+ N_XI12.XI27.NET58_XI12.XI27.MM6_g N_VSS_XI12.XI27.MM6_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI22.MM6 N_XI12.XI22.NET15_XI12.XI22.MM6_d
+ N_XI12.XI22.NET58_XI12.XI22.MM6_g N_VSS_XI12.XI22.MM6_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI21.MM6 N_XI12.XI21.NET15_XI12.XI21.MM6_d
+ N_XI12.XI21.NET58_XI12.XI21.MM6_g N_VSS_XI12.XI21.MM6_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI23.MM6 N_XI12.XI23.NET15_XI12.XI23.MM6_d
+ N_XI12.XI23.NET58_XI12.XI23.MM6_g N_VSS_XI12.XI23.MM6_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI19.MM6 N_XI12.XI19.NET15_XI12.XI19.MM6_d
+ N_XI12.XI19.NET58_XI12.XI19.MM6_g N_VSS_XI12.XI19.MM6_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI20.MM6 N_XI12.XI20.NET15_XI12.XI20.MM6_d
+ N_XI12.XI20.NET58_XI12.XI20.MM6_g N_VSS_XI12.XI20.MM6_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI18.MM6 N_XI12.XI18.NET15_XI12.XI18.MM6_d
+ N_XI12.XI18.NET58_XI12.XI18.MM6_g N_VSS_XI12.XI18.MM6_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI17.MM6 N_XI12.XI17.NET15_XI12.XI17.MM6_d
+ N_XI12.XI17.NET58_XI12.XI17.MM6_g N_VSS_XI12.XI17.MM6_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI0.MM6 N_XI12.XI0.NET15_XI12.XI0.MM6_d N_XI12.XI0.NET58_XI12.XI0.MM6_g
+ N_VSS_XI12.XI0.MM6_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI12.XI30.MM0 N_XI12.XI30.NET54_XI12.XI30.MM0_d
+ N_XI12.XI30.NET15_XI12.XI30.MM0_g N_VSS_XI12.XI30.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI29.MM0 N_XI12.XI29.NET54_XI12.XI29.MM0_d
+ N_XI12.XI29.NET15_XI12.XI29.MM0_g N_VSS_XI12.XI29.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI31.MM0 N_XI12.XI31.NET54_XI12.XI31.MM0_d
+ N_XI12.XI31.NET15_XI12.XI31.MM0_g N_VSS_XI12.XI31.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI28.MM0 N_XI12.XI28.NET54_XI12.XI28.MM0_d
+ N_XI12.XI28.NET15_XI12.XI28.MM0_g N_VSS_XI12.XI28.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI25.MM0 N_XI12.XI25.NET54_XI12.XI25.MM0_d
+ N_XI12.XI25.NET15_XI12.XI25.MM0_g N_VSS_XI12.XI25.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI26.MM0 N_XI12.XI26.NET54_XI12.XI26.MM0_d
+ N_XI12.XI26.NET15_XI12.XI26.MM0_g N_VSS_XI12.XI26.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI24.MM0 N_XI12.XI24.NET54_XI12.XI24.MM0_d
+ N_XI12.XI24.NET15_XI12.XI24.MM0_g N_VSS_XI12.XI24.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI27.MM0 N_XI12.XI27.NET54_XI12.XI27.MM0_d
+ N_XI12.XI27.NET15_XI12.XI27.MM0_g N_VSS_XI12.XI27.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI22.MM0 N_XI12.XI22.NET54_XI12.XI22.MM0_d
+ N_XI12.XI22.NET15_XI12.XI22.MM0_g N_VSS_XI12.XI22.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI21.MM0 N_XI12.XI21.NET54_XI12.XI21.MM0_d
+ N_XI12.XI21.NET15_XI12.XI21.MM0_g N_VSS_XI12.XI21.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI23.MM0 N_XI12.XI23.NET54_XI12.XI23.MM0_d
+ N_XI12.XI23.NET15_XI12.XI23.MM0_g N_VSS_XI12.XI23.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI19.MM0 N_XI12.XI19.NET54_XI12.XI19.MM0_d
+ N_XI12.XI19.NET15_XI12.XI19.MM0_g N_VSS_XI12.XI19.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI20.MM0 N_XI12.XI20.NET54_XI12.XI20.MM0_d
+ N_XI12.XI20.NET15_XI12.XI20.MM0_g N_VSS_XI12.XI20.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI18.MM0 N_XI12.XI18.NET54_XI12.XI18.MM0_d
+ N_XI12.XI18.NET15_XI12.XI18.MM0_g N_VSS_XI12.XI18.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI17.MM0 N_XI12.XI17.NET54_XI12.XI17.MM0_d
+ N_XI12.XI17.NET15_XI12.XI17.MM0_g N_VSS_XI12.XI17.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI0.MM0 N_XI12.XI0.NET54_XI12.XI0.MM0_d N_XI12.XI0.NET15_XI12.XI0.MM0_g
+ N_VSS_XI12.XI0.MM0_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI12.XI30.MM36 N_XI12.XI30.NET58_XI12.XI30.MM36_d
+ N_XI12.XI30.NET35_XI12.XI30.MM36_g N_XI12.XI30.NET54_XI12.XI30.MM36_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI29.MM36 N_XI12.XI29.NET58_XI12.XI29.MM36_d
+ N_XI12.XI29.NET35_XI12.XI29.MM36_g N_XI12.XI29.NET54_XI12.XI29.MM36_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI31.MM36 N_XI12.XI31.NET58_XI12.XI31.MM36_d
+ N_XI12.XI31.NET35_XI12.XI31.MM36_g N_XI12.XI31.NET54_XI12.XI31.MM36_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI28.MM36 N_XI12.XI28.NET58_XI12.XI28.MM36_d
+ N_XI12.XI28.NET35_XI12.XI28.MM36_g N_XI12.XI28.NET54_XI12.XI28.MM36_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI25.MM36 N_XI12.XI25.NET58_XI12.XI25.MM36_d
+ N_XI12.XI25.NET35_XI12.XI25.MM36_g N_XI12.XI25.NET54_XI12.XI25.MM36_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI26.MM36 N_XI12.XI26.NET58_XI12.XI26.MM36_d
+ N_XI12.XI26.NET35_XI12.XI26.MM36_g N_XI12.XI26.NET54_XI12.XI26.MM36_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI24.MM36 N_XI12.XI24.NET58_XI12.XI24.MM36_d
+ N_XI12.XI24.NET35_XI12.XI24.MM36_g N_XI12.XI24.NET54_XI12.XI24.MM36_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI27.MM36 N_XI12.XI27.NET58_XI12.XI27.MM36_d
+ N_XI12.XI27.NET35_XI12.XI27.MM36_g N_XI12.XI27.NET54_XI12.XI27.MM36_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI22.MM36 N_XI12.XI22.NET58_XI12.XI22.MM36_d
+ N_XI12.XI22.NET35_XI12.XI22.MM36_g N_XI12.XI22.NET54_XI12.XI22.MM36_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI21.MM36 N_XI12.XI21.NET58_XI12.XI21.MM36_d
+ N_XI12.XI21.NET35_XI12.XI21.MM36_g N_XI12.XI21.NET54_XI12.XI21.MM36_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI23.MM36 N_XI12.XI23.NET58_XI12.XI23.MM36_d
+ N_XI12.XI23.NET35_XI12.XI23.MM36_g N_XI12.XI23.NET54_XI12.XI23.MM36_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI19.MM36 N_XI12.XI19.NET58_XI12.XI19.MM36_d
+ N_XI12.XI19.NET35_XI12.XI19.MM36_g N_XI12.XI19.NET54_XI12.XI19.MM36_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI20.MM36 N_XI12.XI20.NET58_XI12.XI20.MM36_d
+ N_XI12.XI20.NET35_XI12.XI20.MM36_g N_XI12.XI20.NET54_XI12.XI20.MM36_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI18.MM36 N_XI12.XI18.NET58_XI12.XI18.MM36_d
+ N_XI12.XI18.NET35_XI12.XI18.MM36_g N_XI12.XI18.NET54_XI12.XI18.MM36_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI17.MM36 N_XI12.XI17.NET58_XI12.XI17.MM36_d
+ N_XI12.XI17.NET35_XI12.XI17.MM36_g N_XI12.XI17.NET54_XI12.XI17.MM36_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI0.MM36 N_XI12.XI0.NET58_XI12.XI0.MM36_d N_XI12.XI0.NET35_XI12.XI0.MM36_g
+ N_XI12.XI0.NET54_XI12.XI0.MM36_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI12.XI30.MM38 N_XI12.XI30.NET15_XI12.XI30.MM38_d
+ N_XI12.XI30.NET35_XI12.XI30.MM38_g N_XI12.XI30.NET14_XI12.XI30.MM38_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI29.MM38 N_XI12.XI29.NET15_XI12.XI29.MM38_d
+ N_XI12.XI29.NET35_XI12.XI29.MM38_g N_XI12.XI29.NET14_XI12.XI29.MM38_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI31.MM38 N_XI12.XI31.NET15_XI12.XI31.MM38_d
+ N_XI12.XI31.NET35_XI12.XI31.MM38_g N_XI12.XI31.NET14_XI12.XI31.MM38_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI28.MM38 N_XI12.XI28.NET15_XI12.XI28.MM38_d
+ N_XI12.XI28.NET35_XI12.XI28.MM38_g N_XI12.XI28.NET14_XI12.XI28.MM38_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI25.MM38 N_XI12.XI25.NET15_XI12.XI25.MM38_d
+ N_XI12.XI25.NET35_XI12.XI25.MM38_g N_XI12.XI25.NET14_XI12.XI25.MM38_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI26.MM38 N_XI12.XI26.NET15_XI12.XI26.MM38_d
+ N_XI12.XI26.NET35_XI12.XI26.MM38_g N_XI12.XI26.NET14_XI12.XI26.MM38_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI24.MM38 N_XI12.XI24.NET15_XI12.XI24.MM38_d
+ N_XI12.XI24.NET35_XI12.XI24.MM38_g N_XI12.XI24.NET14_XI12.XI24.MM38_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI27.MM38 N_XI12.XI27.NET15_XI12.XI27.MM38_d
+ N_XI12.XI27.NET35_XI12.XI27.MM38_g N_XI12.XI27.NET14_XI12.XI27.MM38_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI22.MM38 N_XI12.XI22.NET15_XI12.XI22.MM38_d
+ N_XI12.XI22.NET35_XI12.XI22.MM38_g N_XI12.XI22.NET14_XI12.XI22.MM38_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI21.MM38 N_XI12.XI21.NET15_XI12.XI21.MM38_d
+ N_XI12.XI21.NET35_XI12.XI21.MM38_g N_XI12.XI21.NET14_XI12.XI21.MM38_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI23.MM38 N_XI12.XI23.NET15_XI12.XI23.MM38_d
+ N_XI12.XI23.NET35_XI12.XI23.MM38_g N_XI12.XI23.NET14_XI12.XI23.MM38_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI19.MM38 N_XI12.XI19.NET15_XI12.XI19.MM38_d
+ N_XI12.XI19.NET35_XI12.XI19.MM38_g N_XI12.XI19.NET14_XI12.XI19.MM38_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI20.MM38 N_XI12.XI20.NET15_XI12.XI20.MM38_d
+ N_XI12.XI20.NET35_XI12.XI20.MM38_g N_XI12.XI20.NET14_XI12.XI20.MM38_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI18.MM38 N_XI12.XI18.NET15_XI12.XI18.MM38_d
+ N_XI12.XI18.NET35_XI12.XI18.MM38_g N_XI12.XI18.NET14_XI12.XI18.MM38_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI17.MM38 N_XI12.XI17.NET15_XI12.XI17.MM38_d
+ N_XI12.XI17.NET35_XI12.XI17.MM38_g N_XI12.XI17.NET14_XI12.XI17.MM38_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI0.MM38 N_XI12.XI0.NET15_XI12.XI0.MM38_d N_XI12.XI0.NET35_XI12.XI0.MM38_g
+ N_XI12.XI0.NET14_XI12.XI0.MM38_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI12.XI30.MM15 N_MIN15_XI12.XI30.MM15_d N_XI12.XI30.NET14_XI12.XI30.MM15_g
+ N_VSS_XI12.XI30.MM15_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI12.XI29.MM15 N_MIN14_XI12.XI29.MM15_d N_XI12.XI29.NET14_XI12.XI29.MM15_g
+ N_VSS_XI12.XI29.MM15_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI12.XI31.MM15 N_MIN13_XI12.XI31.MM15_d N_XI12.XI31.NET14_XI12.XI31.MM15_g
+ N_VSS_XI12.XI31.MM15_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI12.XI28.MM15 N_MIN12_XI12.XI28.MM15_d N_XI12.XI28.NET14_XI12.XI28.MM15_g
+ N_VSS_XI12.XI28.MM15_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI12.XI25.MM15 N_MIN11_XI12.XI25.MM15_d N_XI12.XI25.NET14_XI12.XI25.MM15_g
+ N_VSS_XI12.XI25.MM15_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI12.XI26.MM15 N_MIN10_XI12.XI26.MM15_d N_XI12.XI26.NET14_XI12.XI26.MM15_g
+ N_VSS_XI12.XI26.MM15_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI12.XI24.MM15 N_MIN9_XI12.XI24.MM15_d N_XI12.XI24.NET14_XI12.XI24.MM15_g
+ N_VSS_XI12.XI24.MM15_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI12.XI27.MM15 N_MIN8_XI12.XI27.MM15_d N_XI12.XI27.NET14_XI12.XI27.MM15_g
+ N_VSS_XI12.XI27.MM15_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI12.XI22.MM15 N_MIN7_XI12.XI22.MM15_d N_XI12.XI22.NET14_XI12.XI22.MM15_g
+ N_VSS_XI12.XI22.MM15_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI12.XI21.MM15 N_MIN6_XI12.XI21.MM15_d N_XI12.XI21.NET14_XI12.XI21.MM15_g
+ N_VSS_XI12.XI21.MM15_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI12.XI23.MM15 N_MIN5_XI12.XI23.MM15_d N_XI12.XI23.NET14_XI12.XI23.MM15_g
+ N_VSS_XI12.XI23.MM15_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI12.XI19.MM15 N_MIN4_XI12.XI19.MM15_d N_XI12.XI19.NET14_XI12.XI19.MM15_g
+ N_VSS_XI12.XI19.MM15_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI12.XI20.MM15 N_MIN3_XI12.XI20.MM15_d N_XI12.XI20.NET14_XI12.XI20.MM15_g
+ N_VSS_XI12.XI20.MM15_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI12.XI18.MM15 N_MIN2_XI12.XI18.MM15_d N_XI12.XI18.NET14_XI12.XI18.MM15_g
+ N_VSS_XI12.XI18.MM15_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI12.XI17.MM15 N_MIN1_XI12.XI17.MM15_d N_XI12.XI17.NET14_XI12.XI17.MM15_g
+ N_VSS_XI12.XI17.MM15_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI12.XI0.MM15 N_MIN0_XI12.XI0.MM15_d N_XI12.XI0.NET14_XI12.XI0.MM15_g
+ N_VSS_XI12.XI0.MM15_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI12.XI30.MM16 N_XI12.BAR_Q16_XI12.XI30.MM16_d N_MIN15_XI12.XI30.MM16_g
+ N_VSS_XI12.XI30.MM16_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI12.XI29.MM16 N_XI12.BAR_Q15_XI12.XI29.MM16_d N_MIN14_XI12.XI29.MM16_g
+ N_VSS_XI12.XI29.MM16_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI12.XI31.MM16 N_XI12.BAR_Q14_XI12.XI31.MM16_d N_MIN13_XI12.XI31.MM16_g
+ N_VSS_XI12.XI31.MM16_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI12.XI28.MM16 N_XI12.BAR_Q13_XI12.XI28.MM16_d N_MIN12_XI12.XI28.MM16_g
+ N_VSS_XI12.XI28.MM16_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI12.XI25.MM16 N_XI12.BAR_Q12_XI12.XI25.MM16_d N_MIN11_XI12.XI25.MM16_g
+ N_VSS_XI12.XI25.MM16_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI12.XI26.MM16 N_XI12.BAR_Q11_XI12.XI26.MM16_d N_MIN10_XI12.XI26.MM16_g
+ N_VSS_XI12.XI26.MM16_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI12.XI24.MM16 N_XI12.BAR_Q10_XI12.XI24.MM16_d N_MIN9_XI12.XI24.MM16_g
+ N_VSS_XI12.XI24.MM16_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI12.XI27.MM16 N_XI12.BAR_Q9_XI12.XI27.MM16_d N_MIN8_XI12.XI27.MM16_g
+ N_VSS_XI12.XI27.MM16_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI12.XI22.MM16 N_XI12.BAR_Q8_XI12.XI22.MM16_d N_MIN7_XI12.XI22.MM16_g
+ N_VSS_XI12.XI22.MM16_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI12.XI21.MM16 N_XI12.BAR_Q7_XI12.XI21.MM16_d N_MIN6_XI12.XI21.MM16_g
+ N_VSS_XI12.XI21.MM16_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI12.XI23.MM16 N_XI12.BAR_Q6_XI12.XI23.MM16_d N_MIN5_XI12.XI23.MM16_g
+ N_VSS_XI12.XI23.MM16_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI12.XI19.MM16 N_XI12.BAR_Q5_XI12.XI19.MM16_d N_MIN4_XI12.XI19.MM16_g
+ N_VSS_XI12.XI19.MM16_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI12.XI20.MM16 N_XI12.BAR_Q4_XI12.XI20.MM16_d N_MIN3_XI12.XI20.MM16_g
+ N_VSS_XI12.XI20.MM16_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI12.XI18.MM16 N_XI12.BAR_Q3_XI12.XI18.MM16_d N_MIN2_XI12.XI18.MM16_g
+ N_VSS_XI12.XI18.MM16_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI12.XI17.MM16 N_XI12.BAR_Q2_XI12.XI17.MM16_d N_MIN1_XI12.XI17.MM16_g
+ N_VSS_XI12.XI17.MM16_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI12.XI0.MM16 N_XI12.BAR_Q1_XI12.XI0.MM16_d N_MIN0_XI12.XI0.MM16_g
+ N_VSS_XI12.XI0.MM16_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI12.XI30.MM40 N_XI12.XI30.NET14_XI12.XI30.MM40_d
+ N_XI12.XI30.CLKB_XI12.XI30.MM40_g N_XI12.BAR_Q16_XI12.XI30.MM40_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI29.MM40 N_XI12.XI29.NET14_XI12.XI29.MM40_d
+ N_XI12.XI29.CLKB_XI12.XI29.MM40_g N_XI12.BAR_Q15_XI12.XI29.MM40_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI31.MM40 N_XI12.XI31.NET14_XI12.XI31.MM40_d
+ N_XI12.XI31.CLKB_XI12.XI31.MM40_g N_XI12.BAR_Q14_XI12.XI31.MM40_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI28.MM40 N_XI12.XI28.NET14_XI12.XI28.MM40_d
+ N_XI12.XI28.CLKB_XI12.XI28.MM40_g N_XI12.BAR_Q13_XI12.XI28.MM40_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI25.MM40 N_XI12.XI25.NET14_XI12.XI25.MM40_d
+ N_XI12.XI25.CLKB_XI12.XI25.MM40_g N_XI12.BAR_Q12_XI12.XI25.MM40_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI26.MM40 N_XI12.XI26.NET14_XI12.XI26.MM40_d
+ N_XI12.XI26.CLKB_XI12.XI26.MM40_g N_XI12.BAR_Q11_XI12.XI26.MM40_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI24.MM40 N_XI12.XI24.NET14_XI12.XI24.MM40_d
+ N_XI12.XI24.CLKB_XI12.XI24.MM40_g N_XI12.BAR_Q10_XI12.XI24.MM40_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI27.MM40 N_XI12.XI27.NET14_XI12.XI27.MM40_d
+ N_XI12.XI27.CLKB_XI12.XI27.MM40_g N_XI12.BAR_Q9_XI12.XI27.MM40_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI22.MM40 N_XI12.XI22.NET14_XI12.XI22.MM40_d
+ N_XI12.XI22.CLKB_XI12.XI22.MM40_g N_XI12.BAR_Q8_XI12.XI22.MM40_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI21.MM40 N_XI12.XI21.NET14_XI12.XI21.MM40_d
+ N_XI12.XI21.CLKB_XI12.XI21.MM40_g N_XI12.BAR_Q7_XI12.XI21.MM40_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI23.MM40 N_XI12.XI23.NET14_XI12.XI23.MM40_d
+ N_XI12.XI23.CLKB_XI12.XI23.MM40_g N_XI12.BAR_Q6_XI12.XI23.MM40_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI19.MM40 N_XI12.XI19.NET14_XI12.XI19.MM40_d
+ N_XI12.XI19.CLKB_XI12.XI19.MM40_g N_XI12.BAR_Q5_XI12.XI19.MM40_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI20.MM40 N_XI12.XI20.NET14_XI12.XI20.MM40_d
+ N_XI12.XI20.CLKB_XI12.XI20.MM40_g N_XI12.BAR_Q4_XI12.XI20.MM40_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI18.MM40 N_XI12.XI18.NET14_XI12.XI18.MM40_d
+ N_XI12.XI18.CLKB_XI12.XI18.MM40_g N_XI12.BAR_Q3_XI12.XI18.MM40_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI17.MM40 N_XI12.XI17.NET14_XI12.XI17.MM40_d
+ N_XI12.XI17.CLKB_XI12.XI17.MM40_g N_XI12.BAR_Q2_XI12.XI17.MM40_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI12.XI0.MM40 N_XI12.XI0.NET14_XI12.XI0.MM40_d N_XI12.XI0.CLKB_XI12.XI0.MM40_g
+ N_XI12.BAR_Q1_XI12.XI0.MM40_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI1.XI134.XI9.MM2 N_XI1.XI134.NET43_XI1.XI134.XI9.MM2_d
+ N_NET628_XI1.XI134.XI9.MM2_g N_VSS_XI1.XI134.XI9.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI1.XI153.XI1.MM2 N_XI1.XI153.XI1.NET036_XI1.XI153.XI1.MM2_d
+ N_NET629_XI1.XI153.XI1.MM2_g N_VSS_XI1.XI153.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.85e-13 AS=2.45e-13
+ PD=7.4e-07 PS=1.48e-06
mXI1.XI154.XI1.MM2 N_XI1.XI154.XI1.NET036_XI1.XI154.XI1.MM2_d
+ N_NET630_XI1.XI154.XI1.MM2_g N_VSS_XI1.XI154.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.85e-13 AS=2.45e-13
+ PD=7.4e-07 PS=1.48e-06
mXI1.XI157.XI1.MM2 N_XI1.XI157.XI1.NET036_XI1.XI157.XI1.MM2_d
+ N_NET631_XI1.XI157.XI1.MM2_g N_VSS_XI1.XI157.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.85e-13 AS=2.45e-13
+ PD=7.4e-07 PS=1.48e-06
mXI1.XI156.XI1.MM2 N_XI1.XI156.XI1.NET036_XI1.XI156.XI1.MM2_d
+ N_NET632_XI1.XI156.XI1.MM2_g N_VSS_XI1.XI156.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.85e-13 AS=2.45e-13
+ PD=7.4e-07 PS=1.48e-06
mXI1.XI155.XI1.MM2 N_XI1.XI155.XI1.NET036_XI1.XI155.XI1.MM2_d
+ N_NET633_XI1.XI155.XI1.MM2_g N_VSS_XI1.XI155.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.85e-13 AS=2.45e-13
+ PD=7.4e-07 PS=1.48e-06
mXI1.XI133.XI1.MM2 N_XI1.XI133.XI1.NET036_XI1.XI133.XI1.MM2_d
+ N_NET634_XI1.XI133.XI1.MM2_g N_VSS_XI1.XI133.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.85e-13 AS=2.45e-13
+ PD=7.4e-07 PS=1.48e-06
mXI1.XI132.XI1.MM2 N_XI1.XI132.XI1.NET036_XI1.XI132.XI1.MM2_d
+ N_NET635_XI1.XI132.XI1.MM2_g N_VSS_XI1.XI132.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.85e-13 AS=2.45e-13
+ PD=7.4e-07 PS=1.48e-06
mXI1.XI131.XI1.MM2 N_XI1.XI131.XI1.NET036_XI1.XI131.XI1.MM2_d
+ N_NET636_XI1.XI131.XI1.MM2_g N_VSS_XI1.XI131.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.85e-13 AS=2.45e-13
+ PD=7.4e-07 PS=1.48e-06
mXI1.XI111.XI1.MM2 N_XI1.XI111.XI1.NET036_XI1.XI111.XI1.MM2_d
+ N_NET637_XI1.XI111.XI1.MM2_g N_VSS_XI1.XI111.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.85e-13 AS=2.45e-13
+ PD=7.4e-07 PS=1.48e-06
mXI1.XI110.XI1.MM2 N_XI1.XI110.XI1.NET036_XI1.XI110.XI1.MM2_d
+ N_NET638_XI1.XI110.XI1.MM2_g N_VSS_XI1.XI110.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.85e-13 AS=2.45e-13
+ PD=7.4e-07 PS=1.48e-06
mXI1.XI103.XI1.MM2 N_XI1.XI103.XI1.NET036_XI1.XI103.XI1.MM2_d
+ N_NET639_XI1.XI103.XI1.MM2_g N_VSS_XI1.XI103.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.85e-13 AS=2.45e-13
+ PD=7.4e-07 PS=1.48e-06
mXI1.XI102.XI1.MM2 N_XI1.XI102.XI1.NET036_XI1.XI102.XI1.MM2_d
+ N_NET640_XI1.XI102.XI1.MM2_g N_VSS_XI1.XI102.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.85e-13 AS=2.45e-13
+ PD=7.4e-07 PS=1.48e-06
mXI1.XI88.XI1.MM2 N_XI1.XI88.XI1.NET036_XI1.XI88.XI1.MM2_d
+ N_NET641_XI1.XI88.XI1.MM2_g N_VSS_XI1.XI88.XI1.MM2_s N_VSS_XI10.XI0.XI0.MM2_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.85e-13 AS=2.45e-13 PD=7.4e-07 PS=1.48e-06
mXI1.XI82.XI1.MM2 N_XI1.XI82.XI1.NET036_XI1.XI82.XI1.MM2_d
+ N_NET642_XI1.XI82.XI1.MM2_g N_VSS_XI1.XI82.XI1.MM2_s N_VSS_XI10.XI0.XI0.MM2_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.85e-13 AS=2.45e-13 PD=7.4e-07 PS=1.48e-06
mXI1.XI10.XI1.MM2 N_XI1.XI10.XI1.NET036_XI1.XI10.XI1.MM2_d
+ N_NET643_XI1.XI10.XI1.MM2_g N_VSS_XI1.XI10.XI1.MM2_s N_VSS_XI10.XI0.XI0.MM2_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.85e-13 AS=2.45e-13 PD=7.4e-07 PS=1.48e-06
mXI1.XI153.XI1.MM0 N_XI1.XI153.NET6_XI1.XI153.XI1.MM0_d
+ N_MAX14_XI1.XI153.XI1.MM0_g N_XI1.XI153.XI1.NET036_XI1.XI153.XI1.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=1.85e-13
+ PD=1.52e-06 PS=7.4e-07
mXI1.XI154.XI1.MM0 N_XI1.XI154.NET6_XI1.XI154.XI1.MM0_d
+ N_MAX13_XI1.XI154.XI1.MM0_g N_XI1.XI154.XI1.NET036_XI1.XI154.XI1.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=1.85e-13
+ PD=1.52e-06 PS=7.4e-07
mXI1.XI157.XI1.MM0 N_XI1.XI157.NET6_XI1.XI157.XI1.MM0_d
+ N_MAX12_XI1.XI157.XI1.MM0_g N_XI1.XI157.XI1.NET036_XI1.XI157.XI1.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=1.85e-13
+ PD=1.52e-06 PS=7.4e-07
mXI1.XI156.XI1.MM0 N_XI1.XI156.NET6_XI1.XI156.XI1.MM0_d
+ N_MAX11_XI1.XI156.XI1.MM0_g N_XI1.XI156.XI1.NET036_XI1.XI156.XI1.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=1.85e-13
+ PD=1.52e-06 PS=7.4e-07
mXI1.XI155.XI1.MM0 N_XI1.XI155.NET6_XI1.XI155.XI1.MM0_d
+ N_MAX10_XI1.XI155.XI1.MM0_g N_XI1.XI155.XI1.NET036_XI1.XI155.XI1.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=1.85e-13
+ PD=1.52e-06 PS=7.4e-07
mXI1.XI133.XI1.MM0 N_XI1.XI133.NET6_XI1.XI133.XI1.MM0_d
+ N_MAX9_XI1.XI133.XI1.MM0_g N_XI1.XI133.XI1.NET036_XI1.XI133.XI1.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=1.85e-13
+ PD=1.52e-06 PS=7.4e-07
mXI1.XI132.XI1.MM0 N_XI1.XI132.NET6_XI1.XI132.XI1.MM0_d
+ N_MAX8_XI1.XI132.XI1.MM0_g N_XI1.XI132.XI1.NET036_XI1.XI132.XI1.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=1.85e-13
+ PD=1.52e-06 PS=7.4e-07
mXI1.XI131.XI1.MM0 N_XI1.XI131.NET6_XI1.XI131.XI1.MM0_d
+ N_MAX7_XI1.XI131.XI1.MM0_g N_XI1.XI131.XI1.NET036_XI1.XI131.XI1.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=1.85e-13
+ PD=1.52e-06 PS=7.4e-07
mXI1.XI111.XI1.MM0 N_XI1.XI111.NET6_XI1.XI111.XI1.MM0_d
+ N_MAX6_XI1.XI111.XI1.MM0_g N_XI1.XI111.XI1.NET036_XI1.XI111.XI1.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=1.85e-13
+ PD=1.52e-06 PS=7.4e-07
mXI1.XI110.XI1.MM0 N_XI1.XI110.NET6_XI1.XI110.XI1.MM0_d
+ N_MAX5_XI1.XI110.XI1.MM0_g N_XI1.XI110.XI1.NET036_XI1.XI110.XI1.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=1.85e-13
+ PD=1.52e-06 PS=7.4e-07
mXI1.XI103.XI1.MM0 N_XI1.XI103.NET6_XI1.XI103.XI1.MM0_d
+ N_MAX4_XI1.XI103.XI1.MM0_g N_XI1.XI103.XI1.NET036_XI1.XI103.XI1.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=1.85e-13
+ PD=1.52e-06 PS=7.4e-07
mXI1.XI102.XI1.MM0 N_XI1.XI102.NET6_XI1.XI102.XI1.MM0_d
+ N_MAX3_XI1.XI102.XI1.MM0_g N_XI1.XI102.XI1.NET036_XI1.XI102.XI1.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=1.85e-13
+ PD=1.52e-06 PS=7.4e-07
mXI1.XI88.XI1.MM0 N_XI1.XI88.NET6_XI1.XI88.XI1.MM0_d N_MAX2_XI1.XI88.XI1.MM0_g
+ N_XI1.XI88.XI1.NET036_XI1.XI88.XI1.MM0_s N_VSS_XI10.XI0.XI0.MM2_b N_18
+ L=1.8e-07 W=5e-07 AD=2.55e-13 AS=1.85e-13 PD=1.52e-06 PS=7.4e-07
mXI1.XI82.XI1.MM0 N_XI1.XI82.NET6_XI1.XI82.XI1.MM0_d N_MAX1_XI1.XI82.XI1.MM0_g
+ N_XI1.XI82.XI1.NET036_XI1.XI82.XI1.MM0_s N_VSS_XI10.XI0.XI0.MM2_b N_18
+ L=1.8e-07 W=5e-07 AD=2.55e-13 AS=1.85e-13 PD=1.52e-06 PS=7.4e-07
mXI1.XI10.XI1.MM0 N_XI1.XI10.NET6_XI1.XI10.XI1.MM0_d N_MAX0_XI1.XI10.XI1.MM0_g
+ N_XI1.XI10.XI1.NET036_XI1.XI10.XI1.MM0_s N_VSS_XI10.XI0.XI0.MM2_b N_18
+ L=1.8e-07 W=5e-07 AD=2.55e-13 AS=1.85e-13 PD=1.52e-06 PS=7.4e-07
mXI1.XI134.MM2 N_XI1.XI134.NET10_XI1.XI134.MM2_d
+ N_XI1.XI134.NET43_XI1.XI134.MM2_g N_VSS_XI1.XI134.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.2375e-13 AS=3.225e-13
+ PD=8.95e-07 PS=1.79e-06
mXI1.XI153.XI0.MM2 N_XI1.G15_XI1.XI153.XI0.MM2_d
+ N_XI1.XI153.NET6_XI1.XI153.XI0.MM2_g N_VSS_XI1.XI153.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI1.XI154.XI0.MM2 N_XI1.G14_XI1.XI154.XI0.MM2_d
+ N_XI1.XI154.NET6_XI1.XI154.XI0.MM2_g N_VSS_XI1.XI154.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI1.XI157.XI0.MM2 N_XI1.G13_XI1.XI157.XI0.MM2_d
+ N_XI1.XI157.NET6_XI1.XI157.XI0.MM2_g N_VSS_XI1.XI157.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI1.XI156.XI0.MM2 N_XI1.G12_XI1.XI156.XI0.MM2_d
+ N_XI1.XI156.NET6_XI1.XI156.XI0.MM2_g N_VSS_XI1.XI156.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI1.XI155.XI0.MM2 N_XI1.G11_XI1.XI155.XI0.MM2_d
+ N_XI1.XI155.NET6_XI1.XI155.XI0.MM2_g N_VSS_XI1.XI155.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI1.XI133.XI0.MM2 N_XI1.G10_XI1.XI133.XI0.MM2_d
+ N_XI1.XI133.NET6_XI1.XI133.XI0.MM2_g N_VSS_XI1.XI133.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI1.XI132.XI0.MM2 N_XI1.G9_XI1.XI132.XI0.MM2_d
+ N_XI1.XI132.NET6_XI1.XI132.XI0.MM2_g N_VSS_XI1.XI132.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI1.XI131.XI0.MM2 N_XI1.G8_XI1.XI131.XI0.MM2_d
+ N_XI1.XI131.NET6_XI1.XI131.XI0.MM2_g N_VSS_XI1.XI131.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI1.XI111.XI0.MM2 N_XI1.G7_XI1.XI111.XI0.MM2_d
+ N_XI1.XI111.NET6_XI1.XI111.XI0.MM2_g N_VSS_XI1.XI111.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI1.XI110.XI0.MM2 N_XI1.G6_XI1.XI110.XI0.MM2_d
+ N_XI1.XI110.NET6_XI1.XI110.XI0.MM2_g N_VSS_XI1.XI110.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI1.XI103.XI0.MM2 N_XI1.G5_XI1.XI103.XI0.MM2_d
+ N_XI1.XI103.NET6_XI1.XI103.XI0.MM2_g N_VSS_XI1.XI103.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI1.XI102.XI0.MM2 N_XI1.G4_XI1.XI102.XI0.MM2_d
+ N_XI1.XI102.NET6_XI1.XI102.XI0.MM2_g N_VSS_XI1.XI102.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI1.XI88.XI0.MM2 N_XI1.G3_XI1.XI88.XI0.MM2_d N_XI1.XI88.NET6_XI1.XI88.XI0.MM2_g
+ N_VSS_XI1.XI88.XI0.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI1.XI82.XI0.MM2 N_XI1.G2_XI1.XI82.XI0.MM2_d N_XI1.XI82.NET6_XI1.XI82.XI0.MM2_g
+ N_VSS_XI1.XI82.XI0.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI1.XI10.XI0.MM2 N_XI1.G1_XI1.XI10.XI0.MM2_d N_XI1.XI10.NET6_XI1.XI10.XI0.MM2_g
+ N_VSS_XI1.XI10.XI0.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI1.XI134.MM7 N_XI1.P16_XI1.XI134.MM7_d N_XI1.XI134.NET39_XI1.XI134.MM7_g
+ N_XI1.XI134.NET10_XI1.XI134.MM7_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=4.75e-13 AS=2.2375e-13 PD=1.9e-06 PS=8.95e-07
mXI1.XI137.XI9.MM2 N_XI1.XI137.NET43_XI1.XI137.XI9.MM2_d
+ N_NET629_XI1.XI137.XI9.MM2_g N_VSS_XI1.XI137.XI9.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI1.XI140.XI9.MM2 N_XI1.XI140.NET43_XI1.XI140.XI9.MM2_d
+ N_NET630_XI1.XI140.XI9.MM2_g N_VSS_XI1.XI140.XI9.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI1.XI149.XI9.MM2 N_XI1.XI149.NET43_XI1.XI149.XI9.MM2_d
+ N_NET631_XI1.XI149.XI9.MM2_g N_VSS_XI1.XI149.XI9.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI1.XI146.XI9.MM2 N_XI1.XI146.NET43_XI1.XI146.XI9.MM2_d
+ N_NET632_XI1.XI146.XI9.MM2_g N_VSS_XI1.XI146.XI9.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI1.XI143.XI9.MM2 N_XI1.XI143.NET43_XI1.XI143.XI9.MM2_d
+ N_NET633_XI1.XI143.XI9.MM2_g N_VSS_XI1.XI143.XI9.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI1.XI128.XI9.MM2 N_XI1.XI128.NET43_XI1.XI128.XI9.MM2_d
+ N_NET634_XI1.XI128.XI9.MM2_g N_VSS_XI1.XI128.XI9.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI1.XI125.XI9.MM2 N_XI1.XI125.NET43_XI1.XI125.XI9.MM2_d
+ N_NET635_XI1.XI125.XI9.MM2_g N_VSS_XI1.XI125.XI9.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI1.XI122.XI9.MM2 N_XI1.XI122.NET43_XI1.XI122.XI9.MM2_d
+ N_NET636_XI1.XI122.XI9.MM2_g N_VSS_XI1.XI122.XI9.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI1.XI114.XI9.MM2 N_XI1.XI114.NET43_XI1.XI114.XI9.MM2_d
+ N_NET637_XI1.XI114.XI9.MM2_g N_VSS_XI1.XI114.XI9.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI1.XI109.XI9.MM2 N_XI1.XI109.NET43_XI1.XI109.XI9.MM2_d
+ N_NET638_XI1.XI109.XI9.MM2_g N_VSS_XI1.XI109.XI9.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI1.XI106.XI9.MM2 N_XI1.XI106.NET43_XI1.XI106.XI9.MM2_d
+ N_NET639_XI1.XI106.XI9.MM2_g N_VSS_XI1.XI106.XI9.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI1.XI101.XI9.MM2 N_XI1.XI101.NET43_XI1.XI101.XI9.MM2_d
+ N_NET640_XI1.XI101.XI9.MM2_g N_VSS_XI1.XI101.XI9.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI1.XI86.XI9.MM2 N_XI1.XI86.NET43_XI1.XI86.XI9.MM2_d
+ N_NET641_XI1.XI86.XI9.MM2_g N_VSS_XI1.XI86.XI9.MM2_s N_VSS_XI10.XI0.XI0.MM2_b
+ N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI1.XI80.XI9.MM2 N_XI1.XI80.NET43_XI1.XI80.XI9.MM2_d
+ N_NET642_XI1.XI80.XI9.MM2_g N_VSS_XI1.XI80.XI9.MM2_s N_VSS_XI10.XI0.XI0.MM2_b
+ N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI1.XI26.XI9.MM2 N_XI1.XI26.NET43_XI1.XI26.XI9.MM2_d
+ N_NET643_XI1.XI26.XI9.MM2_g N_VSS_XI1.XI26.XI9.MM2_s N_VSS_XI10.XI0.XI0.MM2_b
+ N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI1.XI134.MM6 N_XI1.P16_XI1.XI134.MM6_d N_MAX15_XI1.XI134.MM6_g
+ N_XI1.XI134.NET6_XI1.XI134.MM6_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=4.75e-13 AS=1.8125e-13 PD=1.9e-06 PS=7.25e-07
mXI1.XI134.MM0 N_XI1.XI134.NET6_XI1.XI134.MM0_d N_NET628_XI1.XI134.MM0_g
+ N_VSS_XI1.XI134.MM0_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=1.8125e-13 AS=2.575e-13 PD=7.25e-07 PS=1.53e-06
mXI1.XI137.MM2 N_XI1.XI137.NET10_XI1.XI137.MM2_d
+ N_XI1.XI137.NET43_XI1.XI137.MM2_g N_VSS_XI1.XI137.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.2375e-13 AS=3.225e-13
+ PD=8.95e-07 PS=1.79e-06
mXI1.XI140.MM2 N_XI1.XI140.NET10_XI1.XI140.MM2_d
+ N_XI1.XI140.NET43_XI1.XI140.MM2_g N_VSS_XI1.XI140.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.2375e-13 AS=3.225e-13
+ PD=8.95e-07 PS=1.79e-06
mXI1.XI149.MM2 N_XI1.XI149.NET10_XI1.XI149.MM2_d
+ N_XI1.XI149.NET43_XI1.XI149.MM2_g N_VSS_XI1.XI149.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.2375e-13 AS=3.225e-13
+ PD=8.95e-07 PS=1.79e-06
mXI1.XI146.MM2 N_XI1.XI146.NET10_XI1.XI146.MM2_d
+ N_XI1.XI146.NET43_XI1.XI146.MM2_g N_VSS_XI1.XI146.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.2375e-13 AS=3.225e-13
+ PD=8.95e-07 PS=1.79e-06
mXI1.XI143.MM2 N_XI1.XI143.NET10_XI1.XI143.MM2_d
+ N_XI1.XI143.NET43_XI1.XI143.MM2_g N_VSS_XI1.XI143.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.2375e-13 AS=3.225e-13
+ PD=8.95e-07 PS=1.79e-06
mXI1.XI128.MM2 N_XI1.XI128.NET10_XI1.XI128.MM2_d
+ N_XI1.XI128.NET43_XI1.XI128.MM2_g N_VSS_XI1.XI128.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.2375e-13 AS=3.225e-13
+ PD=8.95e-07 PS=1.79e-06
mXI1.XI125.MM2 N_XI1.XI125.NET10_XI1.XI125.MM2_d
+ N_XI1.XI125.NET43_XI1.XI125.MM2_g N_VSS_XI1.XI125.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.2375e-13 AS=3.225e-13
+ PD=8.95e-07 PS=1.79e-06
mXI1.XI122.MM2 N_XI1.XI122.NET10_XI1.XI122.MM2_d
+ N_XI1.XI122.NET43_XI1.XI122.MM2_g N_VSS_XI1.XI122.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.2375e-13 AS=3.225e-13
+ PD=8.95e-07 PS=1.79e-06
mXI1.XI114.MM2 N_XI1.XI114.NET10_XI1.XI114.MM2_d
+ N_XI1.XI114.NET43_XI1.XI114.MM2_g N_VSS_XI1.XI114.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.2375e-13 AS=3.225e-13
+ PD=8.95e-07 PS=1.79e-06
mXI1.XI109.MM2 N_XI1.XI109.NET10_XI1.XI109.MM2_d
+ N_XI1.XI109.NET43_XI1.XI109.MM2_g N_VSS_XI1.XI109.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.2375e-13 AS=3.225e-13
+ PD=8.95e-07 PS=1.79e-06
mXI1.XI106.MM2 N_XI1.XI106.NET10_XI1.XI106.MM2_d
+ N_XI1.XI106.NET43_XI1.XI106.MM2_g N_VSS_XI1.XI106.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.2375e-13 AS=3.225e-13
+ PD=8.95e-07 PS=1.79e-06
mXI1.XI101.MM2 N_XI1.XI101.NET10_XI1.XI101.MM2_d
+ N_XI1.XI101.NET43_XI1.XI101.MM2_g N_VSS_XI1.XI101.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.2375e-13 AS=3.225e-13
+ PD=8.95e-07 PS=1.79e-06
mXI1.XI86.MM2 N_XI1.XI86.NET10_XI1.XI86.MM2_d N_XI1.XI86.NET43_XI1.XI86.MM2_g
+ N_VSS_XI1.XI86.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.2375e-13 AS=3.225e-13 PD=8.95e-07 PS=1.79e-06
mXI1.XI80.MM2 N_XI1.XI80.NET10_XI1.XI80.MM2_d N_XI1.XI80.NET43_XI1.XI80.MM2_g
+ N_VSS_XI1.XI80.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.2375e-13 AS=3.225e-13 PD=8.95e-07 PS=1.79e-06
mXI1.XI26.MM2 N_XI1.XI26.NET10_XI1.XI26.MM2_d N_XI1.XI26.NET43_XI1.XI26.MM2_g
+ N_VSS_XI1.XI26.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.2375e-13 AS=3.225e-13 PD=8.95e-07 PS=1.79e-06
mXI1.XI137.MM7 N_XI1.P15_XI1.XI137.MM7_d N_XI1.XI137.NET39_XI1.XI137.MM7_g
+ N_XI1.XI137.NET10_XI1.XI137.MM7_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=4.75e-13 AS=2.2375e-13 PD=1.9e-06 PS=8.95e-07
mXI1.XI140.MM7 N_XI1.P14_XI1.XI140.MM7_d N_XI1.XI140.NET39_XI1.XI140.MM7_g
+ N_XI1.XI140.NET10_XI1.XI140.MM7_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=4.75e-13 AS=2.2375e-13 PD=1.9e-06 PS=8.95e-07
mXI1.XI149.MM7 N_XI1.P13_XI1.XI149.MM7_d N_XI1.XI149.NET39_XI1.XI149.MM7_g
+ N_XI1.XI149.NET10_XI1.XI149.MM7_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=4.75e-13 AS=2.2375e-13 PD=1.9e-06 PS=8.95e-07
mXI1.XI146.MM7 N_XI1.P12_XI1.XI146.MM7_d N_XI1.XI146.NET39_XI1.XI146.MM7_g
+ N_XI1.XI146.NET10_XI1.XI146.MM7_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=4.75e-13 AS=2.2375e-13 PD=1.9e-06 PS=8.95e-07
mXI1.XI143.MM7 N_XI1.P11_XI1.XI143.MM7_d N_XI1.XI143.NET39_XI1.XI143.MM7_g
+ N_XI1.XI143.NET10_XI1.XI143.MM7_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=4.75e-13 AS=2.2375e-13 PD=1.9e-06 PS=8.95e-07
mXI1.XI128.MM7 N_XI1.P10_XI1.XI128.MM7_d N_XI1.XI128.NET39_XI1.XI128.MM7_g
+ N_XI1.XI128.NET10_XI1.XI128.MM7_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=4.75e-13 AS=2.2375e-13 PD=1.9e-06 PS=8.95e-07
mXI1.XI125.MM7 N_XI1.P9_XI1.XI125.MM7_d N_XI1.XI125.NET39_XI1.XI125.MM7_g
+ N_XI1.XI125.NET10_XI1.XI125.MM7_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=4.75e-13 AS=2.2375e-13 PD=1.9e-06 PS=8.95e-07
mXI1.XI122.MM7 N_XI1.P8_XI1.XI122.MM7_d N_XI1.XI122.NET39_XI1.XI122.MM7_g
+ N_XI1.XI122.NET10_XI1.XI122.MM7_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=4.75e-13 AS=2.2375e-13 PD=1.9e-06 PS=8.95e-07
mXI1.XI114.MM7 N_XI1.P7_XI1.XI114.MM7_d N_XI1.XI114.NET39_XI1.XI114.MM7_g
+ N_XI1.XI114.NET10_XI1.XI114.MM7_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=4.75e-13 AS=2.2375e-13 PD=1.9e-06 PS=8.95e-07
mXI1.XI109.MM7 N_XI1.P6_XI1.XI109.MM7_d N_XI1.XI109.NET39_XI1.XI109.MM7_g
+ N_XI1.XI109.NET10_XI1.XI109.MM7_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=4.75e-13 AS=2.2375e-13 PD=1.9e-06 PS=8.95e-07
mXI1.XI106.MM7 N_XI1.P5_XI1.XI106.MM7_d N_XI1.XI106.NET39_XI1.XI106.MM7_g
+ N_XI1.XI106.NET10_XI1.XI106.MM7_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=4.75e-13 AS=2.2375e-13 PD=1.9e-06 PS=8.95e-07
mXI1.XI101.MM7 N_XI1.P4_XI1.XI101.MM7_d N_XI1.XI101.NET39_XI1.XI101.MM7_g
+ N_XI1.XI101.NET10_XI1.XI101.MM7_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=4.75e-13 AS=2.2375e-13 PD=1.9e-06 PS=8.95e-07
mXI1.XI86.MM7 N_XI1.P3_XI1.XI86.MM7_d N_XI1.XI86.NET39_XI1.XI86.MM7_g
+ N_XI1.XI86.NET10_XI1.XI86.MM7_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=4.75e-13 AS=2.2375e-13 PD=1.9e-06 PS=8.95e-07
mXI1.XI80.MM7 N_XI1.P2_XI1.XI80.MM7_d N_XI1.XI80.NET39_XI1.XI80.MM7_g
+ N_XI1.XI80.NET10_XI1.XI80.MM7_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=4.75e-13 AS=2.2375e-13 PD=1.9e-06 PS=8.95e-07
mXI1.XI26.MM7 N_XI1.P1_XI1.XI26.MM7_d N_XI1.XI26.NET39_XI1.XI26.MM7_g
+ N_XI1.XI26.NET10_XI1.XI26.MM7_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=4.75e-13 AS=2.2375e-13 PD=1.9e-06 PS=8.95e-07
mXI1.XI134.XI4.MM2 N_XI1.XI134.NET39_XI1.XI134.XI4.MM2_d
+ N_MAX15_XI1.XI134.XI4.MM2_g N_VSS_XI1.XI134.XI4.MM2_s N_VSS_XI10.XI0.XI0.MM2_b
+ N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI1.XI137.MM6 N_XI1.P15_XI1.XI137.MM6_d N_MAX14_XI1.XI137.MM6_g
+ N_XI1.XI137.NET6_XI1.XI137.MM6_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=4.75e-13 AS=1.8125e-13 PD=1.9e-06 PS=7.25e-07
mXI1.XI140.MM6 N_XI1.P14_XI1.XI140.MM6_d N_MAX13_XI1.XI140.MM6_g
+ N_XI1.XI140.NET6_XI1.XI140.MM6_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=4.75e-13 AS=1.8125e-13 PD=1.9e-06 PS=7.25e-07
mXI1.XI149.MM6 N_XI1.P13_XI1.XI149.MM6_d N_MAX12_XI1.XI149.MM6_g
+ N_XI1.XI149.NET6_XI1.XI149.MM6_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=4.75e-13 AS=1.8125e-13 PD=1.9e-06 PS=7.25e-07
mXI1.XI146.MM6 N_XI1.P12_XI1.XI146.MM6_d N_MAX11_XI1.XI146.MM6_g
+ N_XI1.XI146.NET6_XI1.XI146.MM6_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=4.75e-13 AS=1.8125e-13 PD=1.9e-06 PS=7.25e-07
mXI1.XI143.MM6 N_XI1.P11_XI1.XI143.MM6_d N_MAX10_XI1.XI143.MM6_g
+ N_XI1.XI143.NET6_XI1.XI143.MM6_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=4.75e-13 AS=1.8125e-13 PD=1.9e-06 PS=7.25e-07
mXI1.XI128.MM6 N_XI1.P10_XI1.XI128.MM6_d N_MAX9_XI1.XI128.MM6_g
+ N_XI1.XI128.NET6_XI1.XI128.MM6_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=4.75e-13 AS=1.8125e-13 PD=1.9e-06 PS=7.25e-07
mXI1.XI125.MM6 N_XI1.P9_XI1.XI125.MM6_d N_MAX8_XI1.XI125.MM6_g
+ N_XI1.XI125.NET6_XI1.XI125.MM6_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=4.75e-13 AS=1.8125e-13 PD=1.9e-06 PS=7.25e-07
mXI1.XI122.MM6 N_XI1.P8_XI1.XI122.MM6_d N_MAX7_XI1.XI122.MM6_g
+ N_XI1.XI122.NET6_XI1.XI122.MM6_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=4.75e-13 AS=1.8125e-13 PD=1.9e-06 PS=7.25e-07
mXI1.XI114.MM6 N_XI1.P7_XI1.XI114.MM6_d N_MAX6_XI1.XI114.MM6_g
+ N_XI1.XI114.NET6_XI1.XI114.MM6_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=4.75e-13 AS=1.8125e-13 PD=1.9e-06 PS=7.25e-07
mXI1.XI109.MM6 N_XI1.P6_XI1.XI109.MM6_d N_MAX5_XI1.XI109.MM6_g
+ N_XI1.XI109.NET6_XI1.XI109.MM6_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=4.75e-13 AS=1.8125e-13 PD=1.9e-06 PS=7.25e-07
mXI1.XI106.MM6 N_XI1.P5_XI1.XI106.MM6_d N_MAX4_XI1.XI106.MM6_g
+ N_XI1.XI106.NET6_XI1.XI106.MM6_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=4.75e-13 AS=1.8125e-13 PD=1.9e-06 PS=7.25e-07
mXI1.XI101.MM6 N_XI1.P4_XI1.XI101.MM6_d N_MAX3_XI1.XI101.MM6_g
+ N_XI1.XI101.NET6_XI1.XI101.MM6_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=4.75e-13 AS=1.8125e-13 PD=1.9e-06 PS=7.25e-07
mXI1.XI86.MM6 N_XI1.P3_XI1.XI86.MM6_d N_MAX2_XI1.XI86.MM6_g
+ N_XI1.XI86.NET6_XI1.XI86.MM6_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=4.75e-13 AS=1.8125e-13 PD=1.9e-06 PS=7.25e-07
mXI1.XI80.MM6 N_XI1.P2_XI1.XI80.MM6_d N_MAX1_XI1.XI80.MM6_g
+ N_XI1.XI80.NET6_XI1.XI80.MM6_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=4.75e-13 AS=1.8125e-13 PD=1.9e-06 PS=7.25e-07
mXI1.XI26.MM6 N_XI1.P1_XI1.XI26.MM6_d N_MAX0_XI1.XI26.MM6_g
+ N_XI1.XI26.NET6_XI1.XI26.MM6_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=4.75e-13 AS=1.8125e-13 PD=1.9e-06 PS=7.25e-07
mXI1.XI137.MM0 N_XI1.XI137.NET6_XI1.XI137.MM0_d N_NET629_XI1.XI137.MM0_g
+ N_VSS_XI1.XI137.MM0_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=1.8125e-13 AS=2.575e-13 PD=7.25e-07 PS=1.53e-06
mXI1.XI140.MM0 N_XI1.XI140.NET6_XI1.XI140.MM0_d N_NET630_XI1.XI140.MM0_g
+ N_VSS_XI1.XI140.MM0_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=1.8125e-13 AS=2.575e-13 PD=7.25e-07 PS=1.53e-06
mXI1.XI149.MM0 N_XI1.XI149.NET6_XI1.XI149.MM0_d N_NET631_XI1.XI149.MM0_g
+ N_VSS_XI1.XI149.MM0_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=1.8125e-13 AS=2.575e-13 PD=7.25e-07 PS=1.53e-06
mXI1.XI146.MM0 N_XI1.XI146.NET6_XI1.XI146.MM0_d N_NET632_XI1.XI146.MM0_g
+ N_VSS_XI1.XI146.MM0_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=1.8125e-13 AS=2.575e-13 PD=7.25e-07 PS=1.53e-06
mXI1.XI143.MM0 N_XI1.XI143.NET6_XI1.XI143.MM0_d N_NET633_XI1.XI143.MM0_g
+ N_VSS_XI1.XI143.MM0_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=1.8125e-13 AS=2.575e-13 PD=7.25e-07 PS=1.53e-06
mXI1.XI128.MM0 N_XI1.XI128.NET6_XI1.XI128.MM0_d N_NET634_XI1.XI128.MM0_g
+ N_VSS_XI1.XI128.MM0_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=1.8125e-13 AS=2.575e-13 PD=7.25e-07 PS=1.53e-06
mXI1.XI125.MM0 N_XI1.XI125.NET6_XI1.XI125.MM0_d N_NET635_XI1.XI125.MM0_g
+ N_VSS_XI1.XI125.MM0_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=1.8125e-13 AS=2.575e-13 PD=7.25e-07 PS=1.53e-06
mXI1.XI122.MM0 N_XI1.XI122.NET6_XI1.XI122.MM0_d N_NET636_XI1.XI122.MM0_g
+ N_VSS_XI1.XI122.MM0_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=1.8125e-13 AS=2.575e-13 PD=7.25e-07 PS=1.53e-06
mXI1.XI114.MM0 N_XI1.XI114.NET6_XI1.XI114.MM0_d N_NET637_XI1.XI114.MM0_g
+ N_VSS_XI1.XI114.MM0_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=1.8125e-13 AS=2.575e-13 PD=7.25e-07 PS=1.53e-06
mXI1.XI109.MM0 N_XI1.XI109.NET6_XI1.XI109.MM0_d N_NET638_XI1.XI109.MM0_g
+ N_VSS_XI1.XI109.MM0_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=1.8125e-13 AS=2.575e-13 PD=7.25e-07 PS=1.53e-06
mXI1.XI106.MM0 N_XI1.XI106.NET6_XI1.XI106.MM0_d N_NET639_XI1.XI106.MM0_g
+ N_VSS_XI1.XI106.MM0_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=1.8125e-13 AS=2.575e-13 PD=7.25e-07 PS=1.53e-06
mXI1.XI101.MM0 N_XI1.XI101.NET6_XI1.XI101.MM0_d N_NET640_XI1.XI101.MM0_g
+ N_VSS_XI1.XI101.MM0_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=1.8125e-13 AS=2.575e-13 PD=7.25e-07 PS=1.53e-06
mXI1.XI86.MM0 N_XI1.XI86.NET6_XI1.XI86.MM0_d N_NET641_XI1.XI86.MM0_g
+ N_VSS_XI1.XI86.MM0_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=1.8125e-13 AS=2.575e-13 PD=7.25e-07 PS=1.53e-06
mXI1.XI80.MM0 N_XI1.XI80.NET6_XI1.XI80.MM0_d N_NET642_XI1.XI80.MM0_g
+ N_VSS_XI1.XI80.MM0_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=1.8125e-13 AS=2.575e-13 PD=7.25e-07 PS=1.53e-06
mXI1.XI26.MM0 N_XI1.XI26.NET6_XI1.XI26.MM0_d N_NET643_XI1.XI26.MM0_g
+ N_VSS_XI1.XI26.MM0_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=1.8125e-13 AS=2.575e-13 PD=7.25e-07 PS=1.53e-06
mXI3.MM2 N_NET01249_XI3.MM2_d N_NET0855_XI3.MM2_g N_VSS_XI3.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=3e-06 AD=1.47e-12 AS=1.47e-12
+ PD=3.98e-06 PS=3.98e-06
mXI1.XI182.XI9.MM2 N_XI1.XI182.NET43_XI1.XI182.XI9.MM2_d
+ N_XI1.P16_XI1.XI182.XI9.MM2_g N_VSS_XI1.XI182.XI9.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI1.XI137.XI4.MM2 N_XI1.XI137.NET39_XI1.XI137.XI4.MM2_d
+ N_MAX14_XI1.XI137.XI4.MM2_g N_VSS_XI1.XI137.XI4.MM2_s N_VSS_XI10.XI0.XI0.MM2_b
+ N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI1.XI140.XI4.MM2 N_XI1.XI140.NET39_XI1.XI140.XI4.MM2_d
+ N_MAX13_XI1.XI140.XI4.MM2_g N_VSS_XI1.XI140.XI4.MM2_s N_VSS_XI10.XI0.XI0.MM2_b
+ N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI1.XI149.XI4.MM2 N_XI1.XI149.NET39_XI1.XI149.XI4.MM2_d
+ N_MAX12_XI1.XI149.XI4.MM2_g N_VSS_XI1.XI149.XI4.MM2_s N_VSS_XI10.XI0.XI0.MM2_b
+ N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI1.XI146.XI4.MM2 N_XI1.XI146.NET39_XI1.XI146.XI4.MM2_d
+ N_MAX11_XI1.XI146.XI4.MM2_g N_VSS_XI1.XI146.XI4.MM2_s N_VSS_XI10.XI0.XI0.MM2_b
+ N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI1.XI143.XI4.MM2 N_XI1.XI143.NET39_XI1.XI143.XI4.MM2_d
+ N_MAX10_XI1.XI143.XI4.MM2_g N_VSS_XI1.XI143.XI4.MM2_s N_VSS_XI10.XI0.XI0.MM2_b
+ N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI1.XI128.XI4.MM2 N_XI1.XI128.NET39_XI1.XI128.XI4.MM2_d
+ N_MAX9_XI1.XI128.XI4.MM2_g N_VSS_XI1.XI128.XI4.MM2_s N_VSS_XI10.XI0.XI0.MM2_b
+ N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI1.XI125.XI4.MM2 N_XI1.XI125.NET39_XI1.XI125.XI4.MM2_d
+ N_MAX8_XI1.XI125.XI4.MM2_g N_VSS_XI1.XI125.XI4.MM2_s N_VSS_XI10.XI0.XI0.MM2_b
+ N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI1.XI122.XI4.MM2 N_XI1.XI122.NET39_XI1.XI122.XI4.MM2_d
+ N_MAX7_XI1.XI122.XI4.MM2_g N_VSS_XI1.XI122.XI4.MM2_s N_VSS_XI10.XI0.XI0.MM2_b
+ N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI1.XI114.XI4.MM2 N_XI1.XI114.NET39_XI1.XI114.XI4.MM2_d
+ N_MAX6_XI1.XI114.XI4.MM2_g N_VSS_XI1.XI114.XI4.MM2_s N_VSS_XI10.XI0.XI0.MM2_b
+ N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI1.XI109.XI4.MM2 N_XI1.XI109.NET39_XI1.XI109.XI4.MM2_d
+ N_MAX5_XI1.XI109.XI4.MM2_g N_VSS_XI1.XI109.XI4.MM2_s N_VSS_XI10.XI0.XI0.MM2_b
+ N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI1.XI106.XI4.MM2 N_XI1.XI106.NET39_XI1.XI106.XI4.MM2_d
+ N_MAX4_XI1.XI106.XI4.MM2_g N_VSS_XI1.XI106.XI4.MM2_s N_VSS_XI10.XI0.XI0.MM2_b
+ N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI1.XI101.XI4.MM2 N_XI1.XI101.NET39_XI1.XI101.XI4.MM2_d
+ N_MAX3_XI1.XI101.XI4.MM2_g N_VSS_XI1.XI101.XI4.MM2_s N_VSS_XI10.XI0.XI0.MM2_b
+ N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI1.XI86.XI4.MM2 N_XI1.XI86.NET39_XI1.XI86.XI4.MM2_d N_MAX2_XI1.XI86.XI4.MM2_g
+ N_VSS_XI1.XI86.XI4.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI1.XI80.XI4.MM2 N_XI1.XI80.NET39_XI1.XI80.XI4.MM2_d N_MAX1_XI1.XI80.XI4.MM2_g
+ N_VSS_XI1.XI80.XI4.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI1.XI26.XI4.MM2 N_XI1.XI26.NET39_XI1.XI26.XI4.MM2_d N_MAX0_XI1.XI26.XI4.MM2_g
+ N_VSS_XI1.XI26.XI4.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI1.XI182.MM2 N_XI1.XI182.NET10_XI1.XI182.MM2_d
+ N_XI1.XI182.NET43_XI1.XI182.MM2_g N_VSS_XI1.XI182.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.2375e-13 AS=3.225e-13
+ PD=8.95e-07 PS=1.79e-06
mXI1.XI168.XI1.XI1.MM0 N_XI1.XI168.XI1.XI1.NET036_XI1.XI168.XI1.XI1.MM0_d
+ N_XI1.NET288_XI1.XI168.XI1.XI1.MM0_g N_VSS_XI1.XI168.XI1.XI1.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.85e-13 AS=2.45e-13
+ PD=7.4e-07 PS=1.48e-06
mXI1.XI167.XI1.XI1.MM0 N_XI1.XI167.XI1.XI1.NET036_XI1.XI167.XI1.XI1.MM0_d
+ N_XI1.NET282_XI1.XI167.XI1.XI1.MM0_g N_VSS_XI1.XI167.XI1.XI1.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.85e-13 AS=2.45e-13
+ PD=7.4e-07 PS=1.48e-06
mXI1.XI166.XI1.XI1.MM0 N_XI1.XI166.XI1.XI1.NET036_XI1.XI166.XI1.XI1.MM0_d
+ N_XI1.NET276_XI1.XI166.XI1.XI1.MM0_g N_VSS_XI1.XI166.XI1.XI1.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.85e-13 AS=2.45e-13
+ PD=7.4e-07 PS=1.48e-06
mXI1.XI165.XI1.XI1.MM0 N_XI1.XI165.XI1.XI1.NET036_XI1.XI165.XI1.XI1.MM0_d
+ N_XI1.NET270_XI1.XI165.XI1.XI1.MM0_g N_VSS_XI1.XI165.XI1.XI1.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.85e-13 AS=2.45e-13
+ PD=7.4e-07 PS=1.48e-06
mXI1.XI159.XI1.XI1.MM0 N_XI1.XI159.XI1.XI1.NET036_XI1.XI159.XI1.XI1.MM0_d
+ N_XI1.NET246_XI1.XI159.XI1.XI1.MM0_g N_VSS_XI1.XI159.XI1.XI1.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.85e-13 AS=2.45e-13
+ PD=7.4e-07 PS=1.48e-06
mXI1.XI160.XI1.XI1.MM0 N_XI1.XI160.XI1.XI1.NET036_XI1.XI160.XI1.XI1.MM0_d
+ N_XI1.NET252_XI1.XI160.XI1.XI1.MM0_g N_VSS_XI1.XI160.XI1.XI1.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.85e-13 AS=2.45e-13
+ PD=7.4e-07 PS=1.48e-06
mXI1.XI161.XI1.XI1.MM0 N_XI1.XI161.XI1.XI1.NET036_XI1.XI161.XI1.XI1.MM0_d
+ N_XI1.NET258_XI1.XI161.XI1.XI1.MM0_g N_VSS_XI1.XI161.XI1.XI1.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.85e-13 AS=2.45e-13
+ PD=7.4e-07 PS=1.48e-06
mXI1.XI162.XI1.XI1.MM0 N_XI1.XI162.XI1.XI1.NET036_XI1.XI162.XI1.XI1.MM0_d
+ N_XI1.NET264_XI1.XI162.XI1.XI1.MM0_g N_VSS_XI1.XI162.XI1.XI1.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.85e-13 AS=2.45e-13
+ PD=7.4e-07 PS=1.48e-06
mXI1.XI121.XI1.XI1.MM0 N_XI1.XI121.XI1.XI1.NET036_XI1.XI121.XI1.XI1.MM0_d
+ N_XI1.NET204_XI1.XI121.XI1.XI1.MM0_g N_VSS_XI1.XI121.XI1.XI1.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.85e-13 AS=2.45e-13
+ PD=7.4e-07 PS=1.48e-06
mXI1.XI120.XI1.XI1.MM0 N_XI1.XI120.XI1.XI1.NET036_XI1.XI120.XI1.XI1.MM0_d
+ N_XI1.NET210_XI1.XI120.XI1.XI1.MM0_g N_VSS_XI1.XI120.XI1.XI1.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.85e-13 AS=2.45e-13
+ PD=7.4e-07 PS=1.48e-06
mXI1.XI119.XI1.XI1.MM0 N_XI1.XI119.XI1.XI1.NET036_XI1.XI119.XI1.XI1.MM0_d
+ N_XI1.NET216_XI1.XI119.XI1.XI1.MM0_g N_VSS_XI1.XI119.XI1.XI1.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.85e-13 AS=2.45e-13
+ PD=7.4e-07 PS=1.48e-06
mXI1.XI118.XI1.XI1.MM0 N_XI1.XI118.XI1.XI1.NET036_XI1.XI118.XI1.XI1.MM0_d
+ N_XI1.NET222_XI1.XI118.XI1.XI1.MM0_g N_VSS_XI1.XI118.XI1.XI1.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.85e-13 AS=2.45e-13
+ PD=7.4e-07 PS=1.48e-06
mXI1.XI91.XI1.XI1.MM0 N_XI1.XI91.XI1.XI1.NET036_XI1.XI91.XI1.XI1.MM0_d
+ N_XI1.NET228_XI1.XI91.XI1.XI1.MM0_g N_VSS_XI1.XI91.XI1.XI1.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.85e-13 AS=2.45e-13
+ PD=7.4e-07 PS=1.48e-06
mXI1.XI90.XI1.XI1.MM0 N_XI1.XI90.XI1.XI1.NET036_XI1.XI90.XI1.XI1.MM0_d
+ N_XI1.NET240_XI1.XI90.XI1.XI1.MM0_g N_VSS_XI1.XI90.XI1.XI1.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.85e-13 AS=2.45e-13
+ PD=7.4e-07 PS=1.48e-06
mXI1.XI89.XI1.XI1.MM0 N_XI1.XI89.XI1.XI1.NET036_XI1.XI89.XI1.XI1.MM0_d
+ N_CIN2_XI1.XI89.XI1.XI1.MM0_g N_VSS_XI1.XI89.XI1.XI1.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.85e-13 AS=2.45e-13
+ PD=7.4e-07 PS=1.48e-06
mXI1.XI182.MM7 N_NET105_XI1.XI182.MM7_d N_XI1.XI182.NET39_XI1.XI182.MM7_g
+ N_XI1.XI182.NET10_XI1.XI182.MM7_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=4.75e-13 AS=2.2375e-13 PD=1.9e-06 PS=8.95e-07
mXI1.XI168.XI1.XI1.MM2 N_XI1.XI168.XI1.NET6_XI1.XI168.XI1.XI1.MM2_d
+ N_XI1.P15_XI1.XI168.XI1.XI1.MM2_g
+ N_XI1.XI168.XI1.XI1.NET036_XI1.XI168.XI1.XI1.MM2_s N_VSS_XI10.XI0.XI0.MM2_b
+ N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=1.85e-13 PD=1.52e-06 PS=7.4e-07
mXI1.XI167.XI1.XI1.MM2 N_XI1.XI167.XI1.NET6_XI1.XI167.XI1.XI1.MM2_d
+ N_XI1.P14_XI1.XI167.XI1.XI1.MM2_g
+ N_XI1.XI167.XI1.XI1.NET036_XI1.XI167.XI1.XI1.MM2_s N_VSS_XI10.XI0.XI0.MM2_b
+ N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=1.85e-13 PD=1.52e-06 PS=7.4e-07
mXI1.XI166.XI1.XI1.MM2 N_XI1.XI166.XI1.NET6_XI1.XI166.XI1.XI1.MM2_d
+ N_XI1.P13_XI1.XI166.XI1.XI1.MM2_g
+ N_XI1.XI166.XI1.XI1.NET036_XI1.XI166.XI1.XI1.MM2_s N_VSS_XI10.XI0.XI0.MM2_b
+ N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=1.85e-13 PD=1.52e-06 PS=7.4e-07
mXI1.XI165.XI1.XI1.MM2 N_XI1.XI165.XI1.NET6_XI1.XI165.XI1.XI1.MM2_d
+ N_XI1.P12_XI1.XI165.XI1.XI1.MM2_g
+ N_XI1.XI165.XI1.XI1.NET036_XI1.XI165.XI1.XI1.MM2_s N_VSS_XI10.XI0.XI0.MM2_b
+ N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=1.85e-13 PD=1.52e-06 PS=7.4e-07
mXI1.XI159.XI1.XI1.MM2 N_XI1.XI159.XI1.NET6_XI1.XI159.XI1.XI1.MM2_d
+ N_XI1.P11_XI1.XI159.XI1.XI1.MM2_g
+ N_XI1.XI159.XI1.XI1.NET036_XI1.XI159.XI1.XI1.MM2_s N_VSS_XI10.XI0.XI0.MM2_b
+ N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=1.85e-13 PD=1.52e-06 PS=7.4e-07
mXI1.XI160.XI1.XI1.MM2 N_XI1.XI160.XI1.NET6_XI1.XI160.XI1.XI1.MM2_d
+ N_XI1.P10_XI1.XI160.XI1.XI1.MM2_g
+ N_XI1.XI160.XI1.XI1.NET036_XI1.XI160.XI1.XI1.MM2_s N_VSS_XI10.XI0.XI0.MM2_b
+ N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=1.85e-13 PD=1.52e-06 PS=7.4e-07
mXI1.XI161.XI1.XI1.MM2 N_XI1.XI161.XI1.NET6_XI1.XI161.XI1.XI1.MM2_d
+ N_XI1.P9_XI1.XI161.XI1.XI1.MM2_g
+ N_XI1.XI161.XI1.XI1.NET036_XI1.XI161.XI1.XI1.MM2_s N_VSS_XI10.XI0.XI0.MM2_b
+ N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=1.85e-13 PD=1.52e-06 PS=7.4e-07
mXI1.XI162.XI1.XI1.MM2 N_XI1.XI162.XI1.NET6_XI1.XI162.XI1.XI1.MM2_d
+ N_XI1.P8_XI1.XI162.XI1.XI1.MM2_g
+ N_XI1.XI162.XI1.XI1.NET036_XI1.XI162.XI1.XI1.MM2_s N_VSS_XI10.XI0.XI0.MM2_b
+ N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=1.85e-13 PD=1.52e-06 PS=7.4e-07
mXI1.XI121.XI1.XI1.MM2 N_XI1.XI121.XI1.NET6_XI1.XI121.XI1.XI1.MM2_d
+ N_XI1.P7_XI1.XI121.XI1.XI1.MM2_g
+ N_XI1.XI121.XI1.XI1.NET036_XI1.XI121.XI1.XI1.MM2_s N_VSS_XI10.XI0.XI0.MM2_b
+ N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=1.85e-13 PD=1.52e-06 PS=7.4e-07
mXI1.XI120.XI1.XI1.MM2 N_XI1.XI120.XI1.NET6_XI1.XI120.XI1.XI1.MM2_d
+ N_XI1.P6_XI1.XI120.XI1.XI1.MM2_g
+ N_XI1.XI120.XI1.XI1.NET036_XI1.XI120.XI1.XI1.MM2_s N_VSS_XI10.XI0.XI0.MM2_b
+ N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=1.85e-13 PD=1.52e-06 PS=7.4e-07
mXI1.XI119.XI1.XI1.MM2 N_XI1.XI119.XI1.NET6_XI1.XI119.XI1.XI1.MM2_d
+ N_XI1.P5_XI1.XI119.XI1.XI1.MM2_g
+ N_XI1.XI119.XI1.XI1.NET036_XI1.XI119.XI1.XI1.MM2_s N_VSS_XI10.XI0.XI0.MM2_b
+ N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=1.85e-13 PD=1.52e-06 PS=7.4e-07
mXI1.XI118.XI1.XI1.MM2 N_XI1.XI118.XI1.NET6_XI1.XI118.XI1.XI1.MM2_d
+ N_XI1.P4_XI1.XI118.XI1.XI1.MM2_g
+ N_XI1.XI118.XI1.XI1.NET036_XI1.XI118.XI1.XI1.MM2_s N_VSS_XI10.XI0.XI0.MM2_b
+ N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=1.85e-13 PD=1.52e-06 PS=7.4e-07
mXI1.XI91.XI1.XI1.MM2 N_XI1.XI91.XI1.NET6_XI1.XI91.XI1.XI1.MM2_d
+ N_XI1.P3_XI1.XI91.XI1.XI1.MM2_g
+ N_XI1.XI91.XI1.XI1.NET036_XI1.XI91.XI1.XI1.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18
+ L=1.8e-07 W=5e-07 AD=2.55e-13 AS=1.85e-13 PD=1.52e-06 PS=7.4e-07
mXI1.XI90.XI1.XI1.MM2 N_XI1.XI90.XI1.NET6_XI1.XI90.XI1.XI1.MM2_d
+ N_XI1.P2_XI1.XI90.XI1.XI1.MM2_g
+ N_XI1.XI90.XI1.XI1.NET036_XI1.XI90.XI1.XI1.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18
+ L=1.8e-07 W=5e-07 AD=2.55e-13 AS=1.85e-13 PD=1.52e-06 PS=7.4e-07
mXI1.XI89.XI1.XI1.MM2 N_XI1.XI89.XI1.NET6_XI1.XI89.XI1.XI1.MM2_d
+ N_XI1.P1_XI1.XI89.XI1.XI1.MM2_g
+ N_XI1.XI89.XI1.XI1.NET036_XI1.XI89.XI1.XI1.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18
+ L=1.8e-07 W=5e-07 AD=2.55e-13 AS=1.85e-13 PD=1.52e-06 PS=7.4e-07
mXI1.XI182.MM6 N_NET105_XI1.XI182.MM6_d N_XI1.NET198_XI1.XI182.MM6_g
+ N_XI1.XI182.NET6_XI1.XI182.MM6_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=4.75e-13 AS=1.8125e-13 PD=1.9e-06 PS=7.25e-07
mXI1.XI168.XI1.XI0.MM2 N_XI1.XI168.NET13_XI1.XI168.XI1.XI0.MM2_d
+ N_XI1.XI168.XI1.NET6_XI1.XI168.XI1.XI0.MM2_g N_VSS_XI1.XI168.XI1.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI1.XI167.XI1.XI0.MM2 N_XI1.XI167.NET13_XI1.XI167.XI1.XI0.MM2_d
+ N_XI1.XI167.XI1.NET6_XI1.XI167.XI1.XI0.MM2_g N_VSS_XI1.XI167.XI1.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI1.XI166.XI1.XI0.MM2 N_XI1.XI166.NET13_XI1.XI166.XI1.XI0.MM2_d
+ N_XI1.XI166.XI1.NET6_XI1.XI166.XI1.XI0.MM2_g N_VSS_XI1.XI166.XI1.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI1.XI165.XI1.XI0.MM2 N_XI1.XI165.NET13_XI1.XI165.XI1.XI0.MM2_d
+ N_XI1.XI165.XI1.NET6_XI1.XI165.XI1.XI0.MM2_g N_VSS_XI1.XI165.XI1.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI1.XI159.XI1.XI0.MM2 N_XI1.XI159.NET13_XI1.XI159.XI1.XI0.MM2_d
+ N_XI1.XI159.XI1.NET6_XI1.XI159.XI1.XI0.MM2_g N_VSS_XI1.XI159.XI1.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI1.XI160.XI1.XI0.MM2 N_XI1.XI160.NET13_XI1.XI160.XI1.XI0.MM2_d
+ N_XI1.XI160.XI1.NET6_XI1.XI160.XI1.XI0.MM2_g N_VSS_XI1.XI160.XI1.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI1.XI161.XI1.XI0.MM2 N_XI1.XI161.NET13_XI1.XI161.XI1.XI0.MM2_d
+ N_XI1.XI161.XI1.NET6_XI1.XI161.XI1.XI0.MM2_g N_VSS_XI1.XI161.XI1.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI1.XI162.XI1.XI0.MM2 N_XI1.XI162.NET13_XI1.XI162.XI1.XI0.MM2_d
+ N_XI1.XI162.XI1.NET6_XI1.XI162.XI1.XI0.MM2_g N_VSS_XI1.XI162.XI1.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI1.XI121.XI1.XI0.MM2 N_XI1.XI121.NET13_XI1.XI121.XI1.XI0.MM2_d
+ N_XI1.XI121.XI1.NET6_XI1.XI121.XI1.XI0.MM2_g N_VSS_XI1.XI121.XI1.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI1.XI120.XI1.XI0.MM2 N_XI1.XI120.NET13_XI1.XI120.XI1.XI0.MM2_d
+ N_XI1.XI120.XI1.NET6_XI1.XI120.XI1.XI0.MM2_g N_VSS_XI1.XI120.XI1.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI1.XI119.XI1.XI0.MM2 N_XI1.XI119.NET13_XI1.XI119.XI1.XI0.MM2_d
+ N_XI1.XI119.XI1.NET6_XI1.XI119.XI1.XI0.MM2_g N_VSS_XI1.XI119.XI1.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI1.XI118.XI1.XI0.MM2 N_XI1.XI118.NET13_XI1.XI118.XI1.XI0.MM2_d
+ N_XI1.XI118.XI1.NET6_XI1.XI118.XI1.XI0.MM2_g N_VSS_XI1.XI118.XI1.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI1.XI91.XI1.XI0.MM2 N_XI1.XI91.NET13_XI1.XI91.XI1.XI0.MM2_d
+ N_XI1.XI91.XI1.NET6_XI1.XI91.XI1.XI0.MM2_g N_VSS_XI1.XI91.XI1.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI1.XI90.XI1.XI0.MM2 N_XI1.XI90.NET13_XI1.XI90.XI1.XI0.MM2_d
+ N_XI1.XI90.XI1.NET6_XI1.XI90.XI1.XI0.MM2_g N_VSS_XI1.XI90.XI1.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI1.XI89.XI1.XI0.MM2 N_XI1.XI89.NET13_XI1.XI89.XI1.XI0.MM2_d
+ N_XI1.XI89.XI1.NET6_XI1.XI89.XI1.XI0.MM2_g N_VSS_XI1.XI89.XI1.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI1.XI182.MM0 N_XI1.XI182.NET6_XI1.XI182.MM0_d N_XI1.P16_XI1.XI182.MM0_g
+ N_VSS_XI1.XI182.MM0_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=1.8125e-13 AS=2.575e-13 PD=7.25e-07 PS=1.53e-06
mXI1.XI168.XI0.XI0.MM0 N_XI1.XI168.XI0.NET12_XI1.XI168.XI0.XI0.MM0_d
+ N_XI1.XI168.NET13_XI1.XI168.XI0.XI0.MM0_g N_VSS_XI1.XI168.XI0.XI0.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.375e-13 AS=2.45e-13
+ PD=5.5e-07 PS=1.48e-06
mXI1.XI167.XI0.XI0.MM0 N_XI1.XI167.XI0.NET12_XI1.XI167.XI0.XI0.MM0_d
+ N_XI1.XI167.NET13_XI1.XI167.XI0.XI0.MM0_g N_VSS_XI1.XI167.XI0.XI0.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.375e-13 AS=2.45e-13
+ PD=5.5e-07 PS=1.48e-06
mXI1.XI166.XI0.XI0.MM0 N_XI1.XI166.XI0.NET12_XI1.XI166.XI0.XI0.MM0_d
+ N_XI1.XI166.NET13_XI1.XI166.XI0.XI0.MM0_g N_VSS_XI1.XI166.XI0.XI0.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.375e-13 AS=2.45e-13
+ PD=5.5e-07 PS=1.48e-06
mXI1.XI165.XI0.XI0.MM0 N_XI1.XI165.XI0.NET12_XI1.XI165.XI0.XI0.MM0_d
+ N_XI1.XI165.NET13_XI1.XI165.XI0.XI0.MM0_g N_VSS_XI1.XI165.XI0.XI0.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.375e-13 AS=2.45e-13
+ PD=5.5e-07 PS=1.48e-06
mXI1.XI159.XI0.XI0.MM0 N_XI1.XI159.XI0.NET12_XI1.XI159.XI0.XI0.MM0_d
+ N_XI1.XI159.NET13_XI1.XI159.XI0.XI0.MM0_g N_VSS_XI1.XI159.XI0.XI0.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.375e-13 AS=2.45e-13
+ PD=5.5e-07 PS=1.48e-06
mXI1.XI160.XI0.XI0.MM0 N_XI1.XI160.XI0.NET12_XI1.XI160.XI0.XI0.MM0_d
+ N_XI1.XI160.NET13_XI1.XI160.XI0.XI0.MM0_g N_VSS_XI1.XI160.XI0.XI0.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.375e-13 AS=2.45e-13
+ PD=5.5e-07 PS=1.48e-06
mXI1.XI161.XI0.XI0.MM0 N_XI1.XI161.XI0.NET12_XI1.XI161.XI0.XI0.MM0_d
+ N_XI1.XI161.NET13_XI1.XI161.XI0.XI0.MM0_g N_VSS_XI1.XI161.XI0.XI0.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.375e-13 AS=2.45e-13
+ PD=5.5e-07 PS=1.48e-06
mXI1.XI162.XI0.XI0.MM0 N_XI1.XI162.XI0.NET12_XI1.XI162.XI0.XI0.MM0_d
+ N_XI1.XI162.NET13_XI1.XI162.XI0.XI0.MM0_g N_VSS_XI1.XI162.XI0.XI0.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.375e-13 AS=2.45e-13
+ PD=5.5e-07 PS=1.48e-06
mXI1.XI121.XI0.XI0.MM0 N_XI1.XI121.XI0.NET12_XI1.XI121.XI0.XI0.MM0_d
+ N_XI1.XI121.NET13_XI1.XI121.XI0.XI0.MM0_g N_VSS_XI1.XI121.XI0.XI0.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.375e-13 AS=2.45e-13
+ PD=5.5e-07 PS=1.48e-06
mXI1.XI120.XI0.XI0.MM0 N_XI1.XI120.XI0.NET12_XI1.XI120.XI0.XI0.MM0_d
+ N_XI1.XI120.NET13_XI1.XI120.XI0.XI0.MM0_g N_VSS_XI1.XI120.XI0.XI0.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.375e-13 AS=2.45e-13
+ PD=5.5e-07 PS=1.48e-06
mXI1.XI119.XI0.XI0.MM0 N_XI1.XI119.XI0.NET12_XI1.XI119.XI0.XI0.MM0_d
+ N_XI1.XI119.NET13_XI1.XI119.XI0.XI0.MM0_g N_VSS_XI1.XI119.XI0.XI0.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.375e-13 AS=2.45e-13
+ PD=5.5e-07 PS=1.48e-06
mXI1.XI118.XI0.XI0.MM0 N_XI1.XI118.XI0.NET12_XI1.XI118.XI0.XI0.MM0_d
+ N_XI1.XI118.NET13_XI1.XI118.XI0.XI0.MM0_g N_VSS_XI1.XI118.XI0.XI0.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.375e-13 AS=2.45e-13
+ PD=5.5e-07 PS=1.48e-06
mXI1.XI91.XI0.XI0.MM0 N_XI1.XI91.XI0.NET12_XI1.XI91.XI0.XI0.MM0_d
+ N_XI1.XI91.NET13_XI1.XI91.XI0.XI0.MM0_g N_VSS_XI1.XI91.XI0.XI0.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.375e-13 AS=2.45e-13
+ PD=5.5e-07 PS=1.48e-06
mXI1.XI90.XI0.XI0.MM0 N_XI1.XI90.XI0.NET12_XI1.XI90.XI0.XI0.MM0_d
+ N_XI1.XI90.NET13_XI1.XI90.XI0.XI0.MM0_g N_VSS_XI1.XI90.XI0.XI0.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.375e-13 AS=2.45e-13
+ PD=5.5e-07 PS=1.48e-06
mXI1.XI89.XI0.XI0.MM0 N_XI1.XI89.XI0.NET12_XI1.XI89.XI0.XI0.MM0_d
+ N_XI1.XI89.NET13_XI1.XI89.XI0.XI0.MM0_g N_VSS_XI1.XI89.XI0.XI0.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.375e-13 AS=2.45e-13
+ PD=5.5e-07 PS=1.48e-06
mXI1.XI182.XI4.MM2 N_XI1.XI182.NET39_XI1.XI182.XI4.MM2_d
+ N_XI1.NET198_XI1.XI182.XI4.MM2_g N_VSS_XI1.XI182.XI4.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI7.MM2 N_NET0855_XI7.MM2_d N_NET105_XI7.MM2_g N_VSS_XI7.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI1.XI168.XI0.XI0.MM2 N_XI1.XI168.XI0.NET12_XI1.XI168.XI0.XI0.MM2_d
+ N_XI1.G15_XI1.XI168.XI0.XI0.MM2_g N_VSS_XI1.XI168.XI0.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.375e-13 AS=2.55e-13
+ PD=5.5e-07 PS=1.52e-06
mXI1.XI167.XI0.XI0.MM2 N_XI1.XI167.XI0.NET12_XI1.XI167.XI0.XI0.MM2_d
+ N_XI1.G14_XI1.XI167.XI0.XI0.MM2_g N_VSS_XI1.XI167.XI0.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.375e-13 AS=2.55e-13
+ PD=5.5e-07 PS=1.52e-06
mXI1.XI166.XI0.XI0.MM2 N_XI1.XI166.XI0.NET12_XI1.XI166.XI0.XI0.MM2_d
+ N_XI1.G13_XI1.XI166.XI0.XI0.MM2_g N_VSS_XI1.XI166.XI0.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.375e-13 AS=2.55e-13
+ PD=5.5e-07 PS=1.52e-06
mXI1.XI165.XI0.XI0.MM2 N_XI1.XI165.XI0.NET12_XI1.XI165.XI0.XI0.MM2_d
+ N_XI1.G12_XI1.XI165.XI0.XI0.MM2_g N_VSS_XI1.XI165.XI0.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.375e-13 AS=2.55e-13
+ PD=5.5e-07 PS=1.52e-06
mXI1.XI159.XI0.XI0.MM2 N_XI1.XI159.XI0.NET12_XI1.XI159.XI0.XI0.MM2_d
+ N_XI1.G11_XI1.XI159.XI0.XI0.MM2_g N_VSS_XI1.XI159.XI0.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.375e-13 AS=2.55e-13
+ PD=5.5e-07 PS=1.52e-06
mXI1.XI160.XI0.XI0.MM2 N_XI1.XI160.XI0.NET12_XI1.XI160.XI0.XI0.MM2_d
+ N_XI1.G10_XI1.XI160.XI0.XI0.MM2_g N_VSS_XI1.XI160.XI0.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.375e-13 AS=2.55e-13
+ PD=5.5e-07 PS=1.52e-06
mXI1.XI161.XI0.XI0.MM2 N_XI1.XI161.XI0.NET12_XI1.XI161.XI0.XI0.MM2_d
+ N_XI1.G9_XI1.XI161.XI0.XI0.MM2_g N_VSS_XI1.XI161.XI0.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.375e-13 AS=2.55e-13
+ PD=5.5e-07 PS=1.52e-06
mXI1.XI162.XI0.XI0.MM2 N_XI1.XI162.XI0.NET12_XI1.XI162.XI0.XI0.MM2_d
+ N_XI1.G8_XI1.XI162.XI0.XI0.MM2_g N_VSS_XI1.XI162.XI0.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.375e-13 AS=2.55e-13
+ PD=5.5e-07 PS=1.52e-06
mXI1.XI121.XI0.XI0.MM2 N_XI1.XI121.XI0.NET12_XI1.XI121.XI0.XI0.MM2_d
+ N_XI1.G7_XI1.XI121.XI0.XI0.MM2_g N_VSS_XI1.XI121.XI0.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.375e-13 AS=2.55e-13
+ PD=5.5e-07 PS=1.52e-06
mXI1.XI120.XI0.XI0.MM2 N_XI1.XI120.XI0.NET12_XI1.XI120.XI0.XI0.MM2_d
+ N_XI1.G6_XI1.XI120.XI0.XI0.MM2_g N_VSS_XI1.XI120.XI0.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.375e-13 AS=2.55e-13
+ PD=5.5e-07 PS=1.52e-06
mXI1.XI119.XI0.XI0.MM2 N_XI1.XI119.XI0.NET12_XI1.XI119.XI0.XI0.MM2_d
+ N_XI1.G5_XI1.XI119.XI0.XI0.MM2_g N_VSS_XI1.XI119.XI0.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.375e-13 AS=2.55e-13
+ PD=5.5e-07 PS=1.52e-06
mXI1.XI118.XI0.XI0.MM2 N_XI1.XI118.XI0.NET12_XI1.XI118.XI0.XI0.MM2_d
+ N_XI1.G4_XI1.XI118.XI0.XI0.MM2_g N_VSS_XI1.XI118.XI0.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.375e-13 AS=2.55e-13
+ PD=5.5e-07 PS=1.52e-06
mXI1.XI91.XI0.XI0.MM2 N_XI1.XI91.XI0.NET12_XI1.XI91.XI0.XI0.MM2_d
+ N_XI1.G3_XI1.XI91.XI0.XI0.MM2_g N_VSS_XI1.XI91.XI0.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.375e-13 AS=2.55e-13
+ PD=5.5e-07 PS=1.52e-06
mXI1.XI90.XI0.XI0.MM2 N_XI1.XI90.XI0.NET12_XI1.XI90.XI0.XI0.MM2_d
+ N_XI1.G2_XI1.XI90.XI0.XI0.MM2_g N_VSS_XI1.XI90.XI0.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.375e-13 AS=2.55e-13
+ PD=5.5e-07 PS=1.52e-06
mXI1.XI89.XI0.XI0.MM2 N_XI1.XI89.XI0.NET12_XI1.XI89.XI0.XI0.MM2_d
+ N_XI1.G1_XI1.XI89.XI0.XI0.MM2_g N_VSS_XI1.XI89.XI0.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.375e-13 AS=2.55e-13
+ PD=5.5e-07 PS=1.52e-06
mXI1.XI168.XI0.XI1.MM2 N_XI1.NET198_XI1.XI168.XI0.XI1.MM2_d
+ N_XI1.XI168.XI0.NET12_XI1.XI168.XI0.XI1.MM2_g N_VSS_XI1.XI168.XI0.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI1.XI167.XI0.XI1.MM2 N_XI1.NET288_XI1.XI167.XI0.XI1.MM2_d
+ N_XI1.XI167.XI0.NET12_XI1.XI167.XI0.XI1.MM2_g N_VSS_XI1.XI167.XI0.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI1.XI166.XI0.XI1.MM2 N_XI1.NET282_XI1.XI166.XI0.XI1.MM2_d
+ N_XI1.XI166.XI0.NET12_XI1.XI166.XI0.XI1.MM2_g N_VSS_XI1.XI166.XI0.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI1.XI165.XI0.XI1.MM2 N_XI1.NET276_XI1.XI165.XI0.XI1.MM2_d
+ N_XI1.XI165.XI0.NET12_XI1.XI165.XI0.XI1.MM2_g N_VSS_XI1.XI165.XI0.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI1.XI159.XI0.XI1.MM2 N_XI1.NET270_XI1.XI159.XI0.XI1.MM2_d
+ N_XI1.XI159.XI0.NET12_XI1.XI159.XI0.XI1.MM2_g N_VSS_XI1.XI159.XI0.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI1.XI160.XI0.XI1.MM2 N_XI1.NET246_XI1.XI160.XI0.XI1.MM2_d
+ N_XI1.XI160.XI0.NET12_XI1.XI160.XI0.XI1.MM2_g N_VSS_XI1.XI160.XI0.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI1.XI161.XI0.XI1.MM2 N_XI1.NET252_XI1.XI161.XI0.XI1.MM2_d
+ N_XI1.XI161.XI0.NET12_XI1.XI161.XI0.XI1.MM2_g N_VSS_XI1.XI161.XI0.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI1.XI162.XI0.XI1.MM2 N_XI1.NET258_XI1.XI162.XI0.XI1.MM2_d
+ N_XI1.XI162.XI0.NET12_XI1.XI162.XI0.XI1.MM2_g N_VSS_XI1.XI162.XI0.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI1.XI121.XI0.XI1.MM2 N_XI1.NET264_XI1.XI121.XI0.XI1.MM2_d
+ N_XI1.XI121.XI0.NET12_XI1.XI121.XI0.XI1.MM2_g N_VSS_XI1.XI121.XI0.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI1.XI120.XI0.XI1.MM2 N_XI1.NET204_XI1.XI120.XI0.XI1.MM2_d
+ N_XI1.XI120.XI0.NET12_XI1.XI120.XI0.XI1.MM2_g N_VSS_XI1.XI120.XI0.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI1.XI119.XI0.XI1.MM2 N_XI1.NET210_XI1.XI119.XI0.XI1.MM2_d
+ N_XI1.XI119.XI0.NET12_XI1.XI119.XI0.XI1.MM2_g N_VSS_XI1.XI119.XI0.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI1.XI118.XI0.XI1.MM2 N_XI1.NET216_XI1.XI118.XI0.XI1.MM2_d
+ N_XI1.XI118.XI0.NET12_XI1.XI118.XI0.XI1.MM2_g N_VSS_XI1.XI118.XI0.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI1.XI91.XI0.XI1.MM2 N_XI1.NET222_XI1.XI91.XI0.XI1.MM2_d
+ N_XI1.XI91.XI0.NET12_XI1.XI91.XI0.XI1.MM2_g N_VSS_XI1.XI91.XI0.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI1.XI90.XI0.XI1.MM2 N_XI1.NET228_XI1.XI90.XI0.XI1.MM2_d
+ N_XI1.XI90.XI0.NET12_XI1.XI90.XI0.XI1.MM2_g N_VSS_XI1.XI90.XI0.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI1.XI89.XI0.XI1.MM2 N_XI1.NET240_XI1.XI89.XI0.XI1.MM2_d
+ N_XI1.XI89.XI0.NET12_XI1.XI89.XI0.XI1.MM2_g N_VSS_XI1.XI89.XI0.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI19.XI18.MM4 N_XI19.XI18.NET7_XI19.XI18.MM4_d N_NET01249_XI19.XI18.MM4_g
+ N_VSS_XI19.XI18.MM4_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI19.XI19.MM4 N_XI19.XI19.NET7_XI19.XI19.MM4_d N_NET01249_XI19.XI19.MM4_g
+ N_VSS_XI19.XI19.MM4_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI19.XI17.MM4 N_XI19.XI17.NET7_XI19.XI17.MM4_d N_NET01249_XI19.XI17.MM4_g
+ N_VSS_XI19.XI17.MM4_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI19.XI16.MM4 N_XI19.XI16.NET7_XI19.XI16.MM4_d N_NET01249_XI19.XI16.MM4_g
+ N_VSS_XI19.XI16.MM4_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI19.XI21.MM4 N_XI19.XI21.NET7_XI19.XI21.MM4_d N_NET01249_XI19.XI21.MM4_g
+ N_VSS_XI19.XI21.MM4_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI19.XI20.MM4 N_XI19.XI20.NET7_XI19.XI20.MM4_d N_NET01249_XI19.XI20.MM4_g
+ N_VSS_XI19.XI20.MM4_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI19.XI22.MM4 N_XI19.XI22.NET7_XI19.XI22.MM4_d N_NET01249_XI19.XI22.MM4_g
+ N_VSS_XI19.XI22.MM4_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI19.XI6.MM4 N_XI19.XI6.NET7_XI19.XI6.MM4_d N_NET01249_XI19.XI6.MM4_g
+ N_VSS_XI19.XI6.MM4_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI19.XI5.MM4 N_XI19.XI5.NET7_XI19.XI5.MM4_d N_NET01249_XI19.XI5.MM4_g
+ N_VSS_XI19.XI5.MM4_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI19.XI7.MM4 N_XI19.XI7.NET7_XI19.XI7.MM4_d N_NET01249_XI19.XI7.MM4_g
+ N_VSS_XI19.XI7.MM4_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI19.XI8.MM4 N_XI19.XI8.NET7_XI19.XI8.MM4_d N_NET01249_XI19.XI8.MM4_g
+ N_VSS_XI19.XI8.MM4_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI19.XI3.MM4 N_XI19.XI3.NET7_XI19.XI3.MM4_d N_NET01249_XI19.XI3.MM4_g
+ N_VSS_XI19.XI3.MM4_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI19.XI4.MM4 N_XI19.XI4.NET7_XI19.XI4.MM4_d N_NET01249_XI19.XI4.MM4_g
+ N_VSS_XI19.XI4.MM4_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI19.XI2.MM4 N_XI19.XI2.NET7_XI19.XI2.MM4_d N_NET01249_XI19.XI2.MM4_g
+ N_VSS_XI19.XI2.MM4_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI19.XI1.MM4 N_XI19.XI1.NET7_XI19.XI1.MM4_d N_NET01249_XI19.XI1.MM4_g
+ N_VSS_XI19.XI1.MM4_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI19.XI0.MM4 N_XI19.XI0.NET7_XI19.XI0.MM4_d N_NET01249_XI19.XI0.MM4_g
+ N_VSS_XI19.XI0.MM4_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI19.XI18.MM3 N_NET241_XI19.XI18.MM3_d N_NET01249_XI19.XI18.MM3_g
+ N_NET559_XI19.XI18.MM3_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=6.05e-13 AS=3.075e-13 PD=2.92e-06 PS=1.23e-06
mXI19.XI19.MM3 N_NET242_XI19.XI19.MM3_d N_NET01249_XI19.XI19.MM3_g
+ N_NET560_XI19.XI19.MM3_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=6.05e-13 AS=3.075e-13 PD=2.92e-06 PS=1.23e-06
mXI19.XI17.MM3 N_NET243_XI19.XI17.MM3_d N_NET01249_XI19.XI17.MM3_g
+ N_NET561_XI19.XI17.MM3_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=6.05e-13 AS=3.075e-13 PD=2.92e-06 PS=1.23e-06
mXI19.XI16.MM3 N_NET244_XI19.XI16.MM3_d N_NET01249_XI19.XI16.MM3_g
+ N_NET562_XI19.XI16.MM3_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=6.05e-13 AS=3.075e-13 PD=2.92e-06 PS=1.23e-06
mXI19.XI21.MM3 N_NET245_XI19.XI21.MM3_d N_NET01249_XI19.XI21.MM3_g
+ N_NET563_XI19.XI21.MM3_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=6.05e-13 AS=3.075e-13 PD=2.92e-06 PS=1.23e-06
mXI19.XI20.MM3 N_NET246_XI19.XI20.MM3_d N_NET01249_XI19.XI20.MM3_g
+ N_NET564_XI19.XI20.MM3_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=6.05e-13 AS=3.075e-13 PD=2.92e-06 PS=1.23e-06
mXI19.XI22.MM3 N_NET247_XI19.XI22.MM3_d N_NET01249_XI19.XI22.MM3_g
+ N_NET565_XI19.XI22.MM3_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=6.05e-13 AS=3.075e-13 PD=2.92e-06 PS=1.23e-06
mXI19.XI6.MM3 N_NET248_XI19.XI6.MM3_d N_NET01249_XI19.XI6.MM3_g
+ N_NET566_XI19.XI6.MM3_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=6.05e-13 AS=3.075e-13 PD=2.92e-06 PS=1.23e-06
mXI19.XI5.MM3 N_NET249_XI19.XI5.MM3_d N_NET01249_XI19.XI5.MM3_g
+ N_NET567_XI19.XI5.MM3_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=6.05e-13 AS=3.075e-13 PD=2.92e-06 PS=1.23e-06
mXI19.XI7.MM3 N_NET250_XI19.XI7.MM3_d N_NET01249_XI19.XI7.MM3_g
+ N_NET568_XI19.XI7.MM3_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=6.05e-13 AS=3.075e-13 PD=2.92e-06 PS=1.23e-06
mXI19.XI8.MM3 N_NET251_XI19.XI8.MM3_d N_NET01249_XI19.XI8.MM3_g
+ N_NET569_XI19.XI8.MM3_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=6.05e-13 AS=3.075e-13 PD=2.92e-06 PS=1.23e-06
mXI19.XI3.MM3 N_NET252_XI19.XI3.MM3_d N_NET01249_XI19.XI3.MM3_g
+ N_NET570_XI19.XI3.MM3_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=6.05e-13 AS=3.075e-13 PD=2.92e-06 PS=1.23e-06
mXI19.XI4.MM3 N_NET253_XI19.XI4.MM3_d N_NET01249_XI19.XI4.MM3_g
+ N_NET571_XI19.XI4.MM3_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=6.05e-13 AS=3.075e-13 PD=2.92e-06 PS=1.23e-06
mXI19.XI2.MM3 N_NET254_XI19.XI2.MM3_d N_NET01249_XI19.XI2.MM3_g
+ N_NET572_XI19.XI2.MM3_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=6.05e-13 AS=3.075e-13 PD=2.92e-06 PS=1.23e-06
mXI19.XI1.MM3 N_NET255_XI19.XI1.MM3_d N_NET01249_XI19.XI1.MM3_g
+ N_NET573_XI19.XI1.MM3_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=6.05e-13 AS=3.075e-13 PD=2.92e-06 PS=1.23e-06
mXI19.XI0.MM3 N_NET256_XI19.XI0.MM3_d N_NET01249_XI19.XI0.MM3_g
+ N_NET574_XI19.XI0.MM3_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=6.05e-13 AS=3.075e-13 PD=2.92e-06 PS=1.23e-06
mXI19.XI18.MM2 N_MAX15_XI19.XI18.MM2_d N_XI19.XI18.NET7_XI19.XI18.MM2_g
+ N_NET559_XI19.XI18.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=3.075e-13 PD=1.48e-06 PS=1.23e-06
mXI19.XI19.MM2 N_MAX14_XI19.XI19.MM2_d N_XI19.XI19.NET7_XI19.XI19.MM2_g
+ N_NET560_XI19.XI19.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=3.075e-13 PD=1.48e-06 PS=1.23e-06
mXI19.XI17.MM2 N_MAX13_XI19.XI17.MM2_d N_XI19.XI17.NET7_XI19.XI17.MM2_g
+ N_NET561_XI19.XI17.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=3.075e-13 PD=1.48e-06 PS=1.23e-06
mXI19.XI16.MM2 N_MAX12_XI19.XI16.MM2_d N_XI19.XI16.NET7_XI19.XI16.MM2_g
+ N_NET562_XI19.XI16.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=3.075e-13 PD=1.48e-06 PS=1.23e-06
mXI19.XI21.MM2 N_MAX11_XI19.XI21.MM2_d N_XI19.XI21.NET7_XI19.XI21.MM2_g
+ N_NET563_XI19.XI21.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=3.075e-13 PD=1.48e-06 PS=1.23e-06
mXI19.XI20.MM2 N_MAX10_XI19.XI20.MM2_d N_XI19.XI20.NET7_XI19.XI20.MM2_g
+ N_NET564_XI19.XI20.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=3.075e-13 PD=1.48e-06 PS=1.23e-06
mXI19.XI22.MM2 N_MAX9_XI19.XI22.MM2_d N_XI19.XI22.NET7_XI19.XI22.MM2_g
+ N_NET565_XI19.XI22.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=3.075e-13 PD=1.48e-06 PS=1.23e-06
mXI19.XI6.MM2 N_MAX8_XI19.XI6.MM2_d N_XI19.XI6.NET7_XI19.XI6.MM2_g
+ N_NET566_XI19.XI6.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=3.075e-13 PD=1.48e-06 PS=1.23e-06
mXI19.XI5.MM2 N_MAX7_XI19.XI5.MM2_d N_XI19.XI5.NET7_XI19.XI5.MM2_g
+ N_NET567_XI19.XI5.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=3.075e-13 PD=1.48e-06 PS=1.23e-06
mXI19.XI7.MM2 N_MAX6_XI19.XI7.MM2_d N_XI19.XI7.NET7_XI19.XI7.MM2_g
+ N_NET568_XI19.XI7.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=3.075e-13 PD=1.48e-06 PS=1.23e-06
mXI19.XI8.MM2 N_MAX5_XI19.XI8.MM2_d N_XI19.XI8.NET7_XI19.XI8.MM2_g
+ N_NET569_XI19.XI8.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=3.075e-13 PD=1.48e-06 PS=1.23e-06
mXI19.XI3.MM2 N_MAX4_XI19.XI3.MM2_d N_XI19.XI3.NET7_XI19.XI3.MM2_g
+ N_NET570_XI19.XI3.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=3.075e-13 PD=1.48e-06 PS=1.23e-06
mXI19.XI4.MM2 N_MAX3_XI19.XI4.MM2_d N_XI19.XI4.NET7_XI19.XI4.MM2_g
+ N_NET571_XI19.XI4.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=3.075e-13 PD=1.48e-06 PS=1.23e-06
mXI19.XI2.MM2 N_MAX2_XI19.XI2.MM2_d N_XI19.XI2.NET7_XI19.XI2.MM2_g
+ N_NET572_XI19.XI2.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=3.075e-13 PD=1.48e-06 PS=1.23e-06
mXI19.XI1.MM2 N_MAX1_XI19.XI1.MM2_d N_XI19.XI1.NET7_XI19.XI1.MM2_g
+ N_NET573_XI19.XI1.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=3.075e-13 PD=1.48e-06 PS=1.23e-06
mXI19.XI0.MM2 N_MAX0_XI19.XI0.MM2_d N_XI19.XI0.NET7_XI19.XI0.MM2_g
+ N_NET574_XI19.XI0.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=3.075e-13 PD=1.48e-06 PS=1.23e-06
mXI14.MM1 N_XI14.NET116_XI14.MM1_d N_NET198_XI14.MM1_g N_VSS_XI14.MM1_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI14.XI16.XI0.MM2 N_XI14.XI16.NET12_XI14.XI16.XI0.MM2_d
+ N_XI14.NET116_XI14.XI16.XI0.MM2_g N_VSS_XI14.XI16.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.875e-13 AS=2.45e-13
+ PD=7.5e-07 PS=1.48e-06
mXI14.XI16.XI0.MM0 N_XI14.XI16.NET12_XI14.XI16.XI0.MM0_d
+ N_NET559_XI14.XI16.XI0.MM0_g N_VSS_XI14.XI16.XI0.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.875e-13 AS=2.55e-13
+ PD=7.5e-07 PS=1.52e-06
mXI14.XI16.XI1.MM2 N_NET382_XI14.XI16.XI1.MM2_d
+ N_XI14.XI16.NET12_XI14.XI16.XI1.MM2_g N_VSS_XI14.XI16.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI14.XI15.XI1.MM2 N_XI14.XI15.XI1.NET036_XI14.XI15.XI1.MM2_d
+ N_NET198_XI14.XI15.XI1.MM2_g N_VSS_XI14.XI15.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.375e-13 AS=2.45e-13
+ PD=5.5e-07 PS=1.48e-06
mXI14.XI15.XI1.MM0 N_XI14.XI15.NET6_XI14.XI15.XI1.MM0_d
+ N_NET560_XI14.XI15.XI1.MM0_g N_XI14.XI15.XI1.NET036_XI14.XI15.XI1.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=1.375e-13
+ PD=1.52e-06 PS=5.5e-07
mXI14.XI15.XI0.MM2 N_NET383_XI14.XI15.XI0.MM2_d
+ N_XI14.XI15.NET6_XI14.XI15.XI0.MM2_g N_VSS_XI14.XI15.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI14.XI14.XI1.MM2 N_XI14.XI14.XI1.NET036_XI14.XI14.XI1.MM2_d
+ N_NET198_XI14.XI14.XI1.MM2_g N_VSS_XI14.XI14.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.375e-13 AS=2.45e-13
+ PD=5.5e-07 PS=1.48e-06
mXI14.XI14.XI1.MM0 N_XI14.XI14.NET6_XI14.XI14.XI1.MM0_d
+ N_NET561_XI14.XI14.XI1.MM0_g N_XI14.XI14.XI1.NET036_XI14.XI14.XI1.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=1.375e-13
+ PD=1.52e-06 PS=5.5e-07
mXI14.XI14.XI0.MM2 N_NET384_XI14.XI14.XI0.MM2_d
+ N_XI14.XI14.NET6_XI14.XI14.XI0.MM2_g N_VSS_XI14.XI14.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI14.XI13.XI1.MM2 N_XI14.XI13.XI1.NET036_XI14.XI13.XI1.MM2_d
+ N_NET198_XI14.XI13.XI1.MM2_g N_VSS_XI14.XI13.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.375e-13 AS=2.45e-13
+ PD=5.5e-07 PS=1.48e-06
mXI14.XI13.XI1.MM0 N_XI14.XI13.NET6_XI14.XI13.XI1.MM0_d
+ N_NET562_XI14.XI13.XI1.MM0_g N_XI14.XI13.XI1.NET036_XI14.XI13.XI1.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=1.375e-13
+ PD=1.52e-06 PS=5.5e-07
mXI14.XI13.XI0.MM2 N_NET385_XI14.XI13.XI0.MM2_d
+ N_XI14.XI13.NET6_XI14.XI13.XI0.MM2_g N_VSS_XI14.XI13.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI14.XI12.XI1.MM2 N_XI14.XI12.XI1.NET036_XI14.XI12.XI1.MM2_d
+ N_NET198_XI14.XI12.XI1.MM2_g N_VSS_XI14.XI12.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.375e-13 AS=2.45e-13
+ PD=5.5e-07 PS=1.48e-06
mXI14.XI12.XI1.MM0 N_XI14.XI12.NET6_XI14.XI12.XI1.MM0_d
+ N_NET563_XI14.XI12.XI1.MM0_g N_XI14.XI12.XI1.NET036_XI14.XI12.XI1.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=1.375e-13
+ PD=1.52e-06 PS=5.5e-07
mXI14.XI12.XI0.MM2 N_NET386_XI14.XI12.XI0.MM2_d
+ N_XI14.XI12.NET6_XI14.XI12.XI0.MM2_g N_VSS_XI14.XI12.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI14.XI11.XI1.MM2 N_XI14.XI11.XI1.NET036_XI14.XI11.XI1.MM2_d
+ N_NET198_XI14.XI11.XI1.MM2_g N_VSS_XI14.XI11.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.375e-13 AS=2.45e-13
+ PD=5.5e-07 PS=1.48e-06
mXI14.XI11.XI1.MM0 N_XI14.XI11.NET6_XI14.XI11.XI1.MM0_d
+ N_NET564_XI14.XI11.XI1.MM0_g N_XI14.XI11.XI1.NET036_XI14.XI11.XI1.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=1.375e-13
+ PD=1.52e-06 PS=5.5e-07
mXI14.XI11.XI0.MM2 N_NET387_XI14.XI11.XI0.MM2_d
+ N_XI14.XI11.NET6_XI14.XI11.XI0.MM2_g N_VSS_XI14.XI11.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI14.XI10.XI1.MM2 N_XI14.XI10.XI1.NET036_XI14.XI10.XI1.MM2_d
+ N_NET198_XI14.XI10.XI1.MM2_g N_VSS_XI14.XI10.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=1.375e-13 AS=2.45e-13
+ PD=5.5e-07 PS=1.48e-06
mXI14.XI10.XI1.MM0 N_XI14.XI10.NET6_XI14.XI10.XI1.MM0_d
+ N_NET565_XI14.XI10.XI1.MM0_g N_XI14.XI10.XI1.NET036_XI14.XI10.XI1.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.55e-13 AS=1.375e-13
+ PD=1.52e-06 PS=5.5e-07
mXI14.XI10.XI0.MM2 N_NET388_XI14.XI10.XI0.MM2_d
+ N_XI14.XI10.NET6_XI14.XI10.XI0.MM2_g N_VSS_XI14.XI10.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI14.XI9.XI1.MM2 N_XI14.XI9.XI1.NET036_XI14.XI9.XI1.MM2_d
+ N_NET198_XI14.XI9.XI1.MM2_g N_VSS_XI14.XI9.XI1.MM2_s N_VSS_XI10.XI0.XI0.MM2_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.375e-13 AS=2.45e-13 PD=5.5e-07 PS=1.48e-06
mXI14.XI9.XI1.MM0 N_XI14.XI9.NET6_XI14.XI9.XI1.MM0_d N_NET566_XI14.XI9.XI1.MM0_g
+ N_XI14.XI9.XI1.NET036_XI14.XI9.XI1.MM0_s N_VSS_XI10.XI0.XI0.MM2_b N_18
+ L=1.8e-07 W=5e-07 AD=2.55e-13 AS=1.375e-13 PD=1.52e-06 PS=5.5e-07
mXI14.XI9.XI0.MM2 N_NET389_XI14.XI9.XI0.MM2_d N_XI14.XI9.NET6_XI14.XI9.XI0.MM2_g
+ N_VSS_XI14.XI9.XI0.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI14.XI8.XI1.MM2 N_XI14.XI8.XI1.NET036_XI14.XI8.XI1.MM2_d
+ N_NET198_XI14.XI8.XI1.MM2_g N_VSS_XI14.XI8.XI1.MM2_s N_VSS_XI10.XI0.XI0.MM2_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.375e-13 AS=2.45e-13 PD=5.5e-07 PS=1.48e-06
mXI14.XI8.XI1.MM0 N_XI14.XI8.NET6_XI14.XI8.XI1.MM0_d N_NET567_XI14.XI8.XI1.MM0_g
+ N_XI14.XI8.XI1.NET036_XI14.XI8.XI1.MM0_s N_VSS_XI10.XI0.XI0.MM2_b N_18
+ L=1.8e-07 W=5e-07 AD=2.55e-13 AS=1.375e-13 PD=1.52e-06 PS=5.5e-07
mXI14.XI8.XI0.MM2 N_NET390_XI14.XI8.XI0.MM2_d N_XI14.XI8.NET6_XI14.XI8.XI0.MM2_g
+ N_VSS_XI14.XI8.XI0.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI14.XI7.XI1.MM2 N_XI14.XI7.XI1.NET036_XI14.XI7.XI1.MM2_d
+ N_NET198_XI14.XI7.XI1.MM2_g N_VSS_XI14.XI7.XI1.MM2_s N_VSS_XI10.XI0.XI0.MM2_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.375e-13 AS=2.45e-13 PD=5.5e-07 PS=1.48e-06
mXI14.XI7.XI1.MM0 N_XI14.XI7.NET6_XI14.XI7.XI1.MM0_d N_NET568_XI14.XI7.XI1.MM0_g
+ N_XI14.XI7.XI1.NET036_XI14.XI7.XI1.MM0_s N_VSS_XI10.XI0.XI0.MM2_b N_18
+ L=1.8e-07 W=5e-07 AD=2.55e-13 AS=1.375e-13 PD=1.52e-06 PS=5.5e-07
mXI14.XI7.XI0.MM2 N_NET391_XI14.XI7.XI0.MM2_d N_XI14.XI7.NET6_XI14.XI7.XI0.MM2_g
+ N_VSS_XI14.XI7.XI0.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI14.XI6.XI1.MM2 N_XI14.XI6.XI1.NET036_XI14.XI6.XI1.MM2_d
+ N_NET198_XI14.XI6.XI1.MM2_g N_VSS_XI14.XI6.XI1.MM2_s N_VSS_XI10.XI0.XI0.MM2_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.375e-13 AS=2.45e-13 PD=5.5e-07 PS=1.48e-06
mXI14.XI6.XI1.MM0 N_XI14.XI6.NET6_XI14.XI6.XI1.MM0_d N_NET569_XI14.XI6.XI1.MM0_g
+ N_XI14.XI6.XI1.NET036_XI14.XI6.XI1.MM0_s N_VSS_XI10.XI0.XI0.MM2_b N_18
+ L=1.8e-07 W=5e-07 AD=2.55e-13 AS=1.375e-13 PD=1.52e-06 PS=5.5e-07
mXI14.XI6.XI0.MM2 N_NET392_XI14.XI6.XI0.MM2_d N_XI14.XI6.NET6_XI14.XI6.XI0.MM2_g
+ N_VSS_XI14.XI6.XI0.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI14.XI5.XI1.MM2 N_XI14.XI5.XI1.NET036_XI14.XI5.XI1.MM2_d
+ N_NET198_XI14.XI5.XI1.MM2_g N_VSS_XI14.XI5.XI1.MM2_s N_VSS_XI10.XI0.XI0.MM2_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.375e-13 AS=2.45e-13 PD=5.5e-07 PS=1.48e-06
mXI14.XI5.XI1.MM0 N_XI14.XI5.NET6_XI14.XI5.XI1.MM0_d N_NET570_XI14.XI5.XI1.MM0_g
+ N_XI14.XI5.XI1.NET036_XI14.XI5.XI1.MM0_s N_VSS_XI10.XI0.XI0.MM2_b N_18
+ L=1.8e-07 W=5e-07 AD=2.55e-13 AS=1.375e-13 PD=1.52e-06 PS=5.5e-07
mXI14.XI5.XI0.MM2 N_NET393_XI14.XI5.XI0.MM2_d N_XI14.XI5.NET6_XI14.XI5.XI0.MM2_g
+ N_VSS_XI14.XI5.XI0.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI14.XI4.XI1.MM2 N_XI14.XI4.XI1.NET036_XI14.XI4.XI1.MM2_d
+ N_NET198_XI14.XI4.XI1.MM2_g N_VSS_XI14.XI4.XI1.MM2_s N_VSS_XI10.XI0.XI0.MM2_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.375e-13 AS=2.45e-13 PD=5.5e-07 PS=1.48e-06
mXI14.XI4.XI1.MM0 N_XI14.XI4.NET6_XI14.XI4.XI1.MM0_d N_NET571_XI14.XI4.XI1.MM0_g
+ N_XI14.XI4.XI1.NET036_XI14.XI4.XI1.MM0_s N_VSS_XI10.XI0.XI0.MM2_b N_18
+ L=1.8e-07 W=5e-07 AD=2.55e-13 AS=1.375e-13 PD=1.52e-06 PS=5.5e-07
mXI14.XI4.XI0.MM2 N_NET394_XI14.XI4.XI0.MM2_d N_XI14.XI4.NET6_XI14.XI4.XI0.MM2_g
+ N_VSS_XI14.XI4.XI0.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI14.XI3.XI1.MM2 N_XI14.XI3.XI1.NET036_XI14.XI3.XI1.MM2_d
+ N_NET198_XI14.XI3.XI1.MM2_g N_VSS_XI14.XI3.XI1.MM2_s N_VSS_XI10.XI0.XI0.MM2_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.375e-13 AS=2.45e-13 PD=5.5e-07 PS=1.48e-06
mXI14.XI3.XI1.MM0 N_XI14.XI3.NET6_XI14.XI3.XI1.MM0_d N_NET572_XI14.XI3.XI1.MM0_g
+ N_XI14.XI3.XI1.NET036_XI14.XI3.XI1.MM0_s N_VSS_XI10.XI0.XI0.MM2_b N_18
+ L=1.8e-07 W=5e-07 AD=2.55e-13 AS=1.375e-13 PD=1.52e-06 PS=5.5e-07
mXI14.XI3.XI0.MM2 N_NET395_XI14.XI3.XI0.MM2_d N_XI14.XI3.NET6_XI14.XI3.XI0.MM2_g
+ N_VSS_XI14.XI3.XI0.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI14.XI2.XI1.MM2 N_XI14.XI2.XI1.NET036_XI14.XI2.XI1.MM2_d
+ N_NET198_XI14.XI2.XI1.MM2_g N_VSS_XI14.XI2.XI1.MM2_s N_VSS_XI10.XI0.XI0.MM2_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.375e-13 AS=2.45e-13 PD=5.5e-07 PS=1.48e-06
mXI14.XI2.XI1.MM0 N_XI14.XI2.NET6_XI14.XI2.XI1.MM0_d N_NET573_XI14.XI2.XI1.MM0_g
+ N_XI14.XI2.XI1.NET036_XI14.XI2.XI1.MM0_s N_VSS_XI10.XI0.XI0.MM2_b N_18
+ L=1.8e-07 W=5e-07 AD=2.55e-13 AS=1.375e-13 PD=1.52e-06 PS=5.5e-07
mXI14.XI2.XI0.MM2 N_NET396_XI14.XI2.XI0.MM2_d N_XI14.XI2.NET6_XI14.XI2.XI0.MM2_g
+ N_VSS_XI14.XI2.XI0.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI14.XI1.XI1.MM2 N_XI14.XI1.XI1.NET036_XI14.XI1.XI1.MM2_d
+ N_NET198_XI14.XI1.XI1.MM2_g N_VSS_XI14.XI1.XI1.MM2_s N_VSS_XI10.XI0.XI0.MM2_b
+ N_18 L=1.8e-07 W=5e-07 AD=1.375e-13 AS=2.45e-13 PD=5.5e-07 PS=1.48e-06
mXI14.XI1.XI1.MM0 N_XI14.XI1.NET6_XI14.XI1.XI1.MM0_d N_NET574_XI14.XI1.XI1.MM0_g
+ N_XI14.XI1.XI1.NET036_XI14.XI1.XI1.MM0_s N_VSS_XI10.XI0.XI0.MM2_b N_18
+ L=1.8e-07 W=5e-07 AD=2.55e-13 AS=1.375e-13 PD=1.52e-06 PS=5.5e-07
mXI14.XI1.XI0.MM2 N_NET397_XI14.XI1.XI0.MM2_d N_XI14.XI1.NET6_XI14.XI1.XI0.MM2_g
+ N_VSS_XI14.XI1.XI0.MM2_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI13.XI30.XI0.MM2 N_XI13.XI30.NET0180_XI13.XI30.XI0.MM2_d
+ N_NET222_XI13.XI30.XI0.MM2_g N_VSS_XI13.XI30.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI29.XI0.MM2 N_XI13.XI29.NET0180_XI13.XI29.XI0.MM2_d
+ N_NET222_XI13.XI29.XI0.MM2_g N_VSS_XI13.XI29.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI31.XI0.MM2 N_XI13.XI31.NET0180_XI13.XI31.XI0.MM2_d
+ N_NET222_XI13.XI31.XI0.MM2_g N_VSS_XI13.XI31.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI28.XI0.MM2 N_XI13.XI28.NET0180_XI13.XI28.XI0.MM2_d
+ N_NET222_XI13.XI28.XI0.MM2_g N_VSS_XI13.XI28.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI25.XI0.MM2 N_XI13.XI25.NET0180_XI13.XI25.XI0.MM2_d
+ N_NET222_XI13.XI25.XI0.MM2_g N_VSS_XI13.XI25.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI26.XI0.MM2 N_XI13.XI26.NET0180_XI13.XI26.XI0.MM2_d
+ N_NET222_XI13.XI26.XI0.MM2_g N_VSS_XI13.XI26.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI24.XI0.MM2 N_XI13.XI24.NET0180_XI13.XI24.XI0.MM2_d
+ N_NET222_XI13.XI24.XI0.MM2_g N_VSS_XI13.XI24.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI27.XI0.MM2 N_XI13.XI27.NET0180_XI13.XI27.XI0.MM2_d
+ N_NET222_XI13.XI27.XI0.MM2_g N_VSS_XI13.XI27.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI22.XI0.MM2 N_XI13.XI22.NET0180_XI13.XI22.XI0.MM2_d
+ N_NET222_XI13.XI22.XI0.MM2_g N_VSS_XI13.XI22.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI21.XI0.MM2 N_XI13.XI21.NET0180_XI13.XI21.XI0.MM2_d
+ N_NET222_XI13.XI21.XI0.MM2_g N_VSS_XI13.XI21.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI23.XI0.MM2 N_XI13.XI23.NET0180_XI13.XI23.XI0.MM2_d
+ N_NET222_XI13.XI23.XI0.MM2_g N_VSS_XI13.XI23.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI19.XI0.MM2 N_XI13.XI19.NET0180_XI13.XI19.XI0.MM2_d
+ N_NET222_XI13.XI19.XI0.MM2_g N_VSS_XI13.XI19.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI20.XI0.MM2 N_XI13.XI20.NET0180_XI13.XI20.XI0.MM2_d
+ N_NET222_XI13.XI20.XI0.MM2_g N_VSS_XI13.XI20.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI18.XI0.MM2 N_XI13.XI18.NET0180_XI13.XI18.XI0.MM2_d
+ N_NET222_XI13.XI18.XI0.MM2_g N_VSS_XI13.XI18.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI17.XI0.MM2 N_XI13.XI17.NET0180_XI13.XI17.XI0.MM2_d
+ N_NET222_XI13.XI17.XI0.MM2_g N_VSS_XI13.XI17.XI0.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI0.XI0.MM2 N_XI13.XI0.NET0180_XI13.XI0.XI0.MM2_d
+ N_NET222_XI13.XI0.XI0.MM2_g N_VSS_XI13.XI0.XI0.MM2_s N_VSS_XI10.XI0.XI0.MM2_b
+ N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI13.XI30.XI1.MM2 N_XI13.XI30.NET35_XI13.XI30.XI1.MM2_d
+ N_XI13.XI30.NET0180_XI13.XI30.XI1.MM2_g N_VSS_XI13.XI30.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI29.XI1.MM2 N_XI13.XI29.NET35_XI13.XI29.XI1.MM2_d
+ N_XI13.XI29.NET0180_XI13.XI29.XI1.MM2_g N_VSS_XI13.XI29.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI31.XI1.MM2 N_XI13.XI31.NET35_XI13.XI31.XI1.MM2_d
+ N_XI13.XI31.NET0180_XI13.XI31.XI1.MM2_g N_VSS_XI13.XI31.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI28.XI1.MM2 N_XI13.XI28.NET35_XI13.XI28.XI1.MM2_d
+ N_XI13.XI28.NET0180_XI13.XI28.XI1.MM2_g N_VSS_XI13.XI28.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI25.XI1.MM2 N_XI13.XI25.NET35_XI13.XI25.XI1.MM2_d
+ N_XI13.XI25.NET0180_XI13.XI25.XI1.MM2_g N_VSS_XI13.XI25.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI26.XI1.MM2 N_XI13.XI26.NET35_XI13.XI26.XI1.MM2_d
+ N_XI13.XI26.NET0180_XI13.XI26.XI1.MM2_g N_VSS_XI13.XI26.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI24.XI1.MM2 N_XI13.XI24.NET35_XI13.XI24.XI1.MM2_d
+ N_XI13.XI24.NET0180_XI13.XI24.XI1.MM2_g N_VSS_XI13.XI24.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI27.XI1.MM2 N_XI13.XI27.NET35_XI13.XI27.XI1.MM2_d
+ N_XI13.XI27.NET0180_XI13.XI27.XI1.MM2_g N_VSS_XI13.XI27.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI22.XI1.MM2 N_XI13.XI22.NET35_XI13.XI22.XI1.MM2_d
+ N_XI13.XI22.NET0180_XI13.XI22.XI1.MM2_g N_VSS_XI13.XI22.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI21.XI1.MM2 N_XI13.XI21.NET35_XI13.XI21.XI1.MM2_d
+ N_XI13.XI21.NET0180_XI13.XI21.XI1.MM2_g N_VSS_XI13.XI21.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI23.XI1.MM2 N_XI13.XI23.NET35_XI13.XI23.XI1.MM2_d
+ N_XI13.XI23.NET0180_XI13.XI23.XI1.MM2_g N_VSS_XI13.XI23.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI19.XI1.MM2 N_XI13.XI19.NET35_XI13.XI19.XI1.MM2_d
+ N_XI13.XI19.NET0180_XI13.XI19.XI1.MM2_g N_VSS_XI13.XI19.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI20.XI1.MM2 N_XI13.XI20.NET35_XI13.XI20.XI1.MM2_d
+ N_XI13.XI20.NET0180_XI13.XI20.XI1.MM2_g N_VSS_XI13.XI20.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI18.XI1.MM2 N_XI13.XI18.NET35_XI13.XI18.XI1.MM2_d
+ N_XI13.XI18.NET0180_XI13.XI18.XI1.MM2_g N_VSS_XI13.XI18.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI17.XI1.MM2 N_XI13.XI17.NET35_XI13.XI17.XI1.MM2_d
+ N_XI13.XI17.NET0180_XI13.XI17.XI1.MM2_g N_VSS_XI13.XI17.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI0.XI1.MM2 N_XI13.XI0.NET35_XI13.XI0.XI1.MM2_d
+ N_XI13.XI0.NET0180_XI13.XI0.XI1.MM2_g N_VSS_XI13.XI0.XI1.MM2_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI30.MM26 N_XI13.XI30.CLKB_XI13.XI30.MM26_d
+ N_XI13.XI30.NET35_XI13.XI30.MM26_g N_VSS_XI13.XI30.MM26_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI29.MM26 N_XI13.XI29.CLKB_XI13.XI29.MM26_d
+ N_XI13.XI29.NET35_XI13.XI29.MM26_g N_VSS_XI13.XI29.MM26_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI31.MM26 N_XI13.XI31.CLKB_XI13.XI31.MM26_d
+ N_XI13.XI31.NET35_XI13.XI31.MM26_g N_VSS_XI13.XI31.MM26_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI28.MM26 N_XI13.XI28.CLKB_XI13.XI28.MM26_d
+ N_XI13.XI28.NET35_XI13.XI28.MM26_g N_VSS_XI13.XI28.MM26_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI25.MM26 N_XI13.XI25.CLKB_XI13.XI25.MM26_d
+ N_XI13.XI25.NET35_XI13.XI25.MM26_g N_VSS_XI13.XI25.MM26_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI26.MM26 N_XI13.XI26.CLKB_XI13.XI26.MM26_d
+ N_XI13.XI26.NET35_XI13.XI26.MM26_g N_VSS_XI13.XI26.MM26_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI24.MM26 N_XI13.XI24.CLKB_XI13.XI24.MM26_d
+ N_XI13.XI24.NET35_XI13.XI24.MM26_g N_VSS_XI13.XI24.MM26_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI27.MM26 N_XI13.XI27.CLKB_XI13.XI27.MM26_d
+ N_XI13.XI27.NET35_XI13.XI27.MM26_g N_VSS_XI13.XI27.MM26_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI22.MM26 N_XI13.XI22.CLKB_XI13.XI22.MM26_d
+ N_XI13.XI22.NET35_XI13.XI22.MM26_g N_VSS_XI13.XI22.MM26_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI21.MM26 N_XI13.XI21.CLKB_XI13.XI21.MM26_d
+ N_XI13.XI21.NET35_XI13.XI21.MM26_g N_VSS_XI13.XI21.MM26_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI23.MM26 N_XI13.XI23.CLKB_XI13.XI23.MM26_d
+ N_XI13.XI23.NET35_XI13.XI23.MM26_g N_VSS_XI13.XI23.MM26_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI19.MM26 N_XI13.XI19.CLKB_XI13.XI19.MM26_d
+ N_XI13.XI19.NET35_XI13.XI19.MM26_g N_VSS_XI13.XI19.MM26_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI20.MM26 N_XI13.XI20.CLKB_XI13.XI20.MM26_d
+ N_XI13.XI20.NET35_XI13.XI20.MM26_g N_VSS_XI13.XI20.MM26_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI18.MM26 N_XI13.XI18.CLKB_XI13.XI18.MM26_d
+ N_XI13.XI18.NET35_XI13.XI18.MM26_g N_VSS_XI13.XI18.MM26_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI17.MM26 N_XI13.XI17.CLKB_XI13.XI17.MM26_d
+ N_XI13.XI17.NET35_XI13.XI17.MM26_g N_VSS_XI13.XI17.MM26_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI0.MM26 N_XI13.XI0.CLKB_XI13.XI0.MM26_d N_XI13.XI0.NET35_XI13.XI0.MM26_g
+ N_VSS_XI13.XI0.MM26_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI13.XI30.MM19 N_XI13.XI30.NET27_XI13.XI30.MM19_d N_NET382_XI13.XI30.MM19_g
+ N_VSS_XI13.XI30.MM19_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI13.XI29.MM19 N_XI13.XI29.NET27_XI13.XI29.MM19_d N_NET383_XI13.XI29.MM19_g
+ N_VSS_XI13.XI29.MM19_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI13.XI31.MM19 N_XI13.XI31.NET27_XI13.XI31.MM19_d N_NET384_XI13.XI31.MM19_g
+ N_VSS_XI13.XI31.MM19_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI13.XI28.MM19 N_XI13.XI28.NET27_XI13.XI28.MM19_d N_NET385_XI13.XI28.MM19_g
+ N_VSS_XI13.XI28.MM19_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI13.XI25.MM19 N_XI13.XI25.NET27_XI13.XI25.MM19_d N_NET386_XI13.XI25.MM19_g
+ N_VSS_XI13.XI25.MM19_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI13.XI26.MM19 N_XI13.XI26.NET27_XI13.XI26.MM19_d N_NET387_XI13.XI26.MM19_g
+ N_VSS_XI13.XI26.MM19_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI13.XI24.MM19 N_XI13.XI24.NET27_XI13.XI24.MM19_d N_NET388_XI13.XI24.MM19_g
+ N_VSS_XI13.XI24.MM19_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI13.XI27.MM19 N_XI13.XI27.NET27_XI13.XI27.MM19_d N_NET389_XI13.XI27.MM19_g
+ N_VSS_XI13.XI27.MM19_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI13.XI22.MM19 N_XI13.XI22.NET27_XI13.XI22.MM19_d N_NET390_XI13.XI22.MM19_g
+ N_VSS_XI13.XI22.MM19_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI13.XI21.MM19 N_XI13.XI21.NET27_XI13.XI21.MM19_d N_NET391_XI13.XI21.MM19_g
+ N_VSS_XI13.XI21.MM19_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI13.XI23.MM19 N_XI13.XI23.NET27_XI13.XI23.MM19_d N_NET392_XI13.XI23.MM19_g
+ N_VSS_XI13.XI23.MM19_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI13.XI19.MM19 N_XI13.XI19.NET27_XI13.XI19.MM19_d N_NET393_XI13.XI19.MM19_g
+ N_VSS_XI13.XI19.MM19_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI13.XI20.MM19 N_XI13.XI20.NET27_XI13.XI20.MM19_d N_NET394_XI13.XI20.MM19_g
+ N_VSS_XI13.XI20.MM19_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI13.XI18.MM19 N_XI13.XI18.NET27_XI13.XI18.MM19_d N_NET395_XI13.XI18.MM19_g
+ N_VSS_XI13.XI18.MM19_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI13.XI17.MM19 N_XI13.XI17.NET27_XI13.XI17.MM19_d N_NET396_XI13.XI17.MM19_g
+ N_VSS_XI13.XI17.MM19_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI13.XI0.MM19 N_XI13.XI0.NET27_XI13.XI0.MM19_d N_NET397_XI13.XI0.MM19_g
+ N_VSS_XI13.XI0.MM19_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI13.XI30.MM18 N_XI13.XI30.NET31_XI13.XI30.MM18_d
+ N_XI13.XI30.NET27_XI13.XI30.MM18_g N_VSS_XI13.XI30.MM18_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI29.MM18 N_XI13.XI29.NET31_XI13.XI29.MM18_d
+ N_XI13.XI29.NET27_XI13.XI29.MM18_g N_VSS_XI13.XI29.MM18_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI31.MM18 N_XI13.XI31.NET31_XI13.XI31.MM18_d
+ N_XI13.XI31.NET27_XI13.XI31.MM18_g N_VSS_XI13.XI31.MM18_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI28.MM18 N_XI13.XI28.NET31_XI13.XI28.MM18_d
+ N_XI13.XI28.NET27_XI13.XI28.MM18_g N_VSS_XI13.XI28.MM18_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI25.MM18 N_XI13.XI25.NET31_XI13.XI25.MM18_d
+ N_XI13.XI25.NET27_XI13.XI25.MM18_g N_VSS_XI13.XI25.MM18_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI26.MM18 N_XI13.XI26.NET31_XI13.XI26.MM18_d
+ N_XI13.XI26.NET27_XI13.XI26.MM18_g N_VSS_XI13.XI26.MM18_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI24.MM18 N_XI13.XI24.NET31_XI13.XI24.MM18_d
+ N_XI13.XI24.NET27_XI13.XI24.MM18_g N_VSS_XI13.XI24.MM18_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI27.MM18 N_XI13.XI27.NET31_XI13.XI27.MM18_d
+ N_XI13.XI27.NET27_XI13.XI27.MM18_g N_VSS_XI13.XI27.MM18_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI22.MM18 N_XI13.XI22.NET31_XI13.XI22.MM18_d
+ N_XI13.XI22.NET27_XI13.XI22.MM18_g N_VSS_XI13.XI22.MM18_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI21.MM18 N_XI13.XI21.NET31_XI13.XI21.MM18_d
+ N_XI13.XI21.NET27_XI13.XI21.MM18_g N_VSS_XI13.XI21.MM18_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI23.MM18 N_XI13.XI23.NET31_XI13.XI23.MM18_d
+ N_XI13.XI23.NET27_XI13.XI23.MM18_g N_VSS_XI13.XI23.MM18_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI19.MM18 N_XI13.XI19.NET31_XI13.XI19.MM18_d
+ N_XI13.XI19.NET27_XI13.XI19.MM18_g N_VSS_XI13.XI19.MM18_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI20.MM18 N_XI13.XI20.NET31_XI13.XI20.MM18_d
+ N_XI13.XI20.NET27_XI13.XI20.MM18_g N_VSS_XI13.XI20.MM18_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI18.MM18 N_XI13.XI18.NET31_XI13.XI18.MM18_d
+ N_XI13.XI18.NET27_XI13.XI18.MM18_g N_VSS_XI13.XI18.MM18_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI17.MM18 N_XI13.XI17.NET31_XI13.XI17.MM18_d
+ N_XI13.XI17.NET27_XI13.XI17.MM18_g N_VSS_XI13.XI17.MM18_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI0.MM18 N_XI13.XI0.NET31_XI13.XI0.MM18_d N_XI13.XI0.NET27_XI13.XI0.MM18_g
+ N_VSS_XI13.XI0.MM18_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI13.XI30.MM28 N_XI13.XI30.NET31_XI13.XI30.MM28_d
+ N_XI13.XI30.CLKB_XI13.XI30.MM28_g N_XI13.XI30.NET58_XI13.XI30.MM28_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI29.MM28 N_XI13.XI29.NET31_XI13.XI29.MM28_d
+ N_XI13.XI29.CLKB_XI13.XI29.MM28_g N_XI13.XI29.NET58_XI13.XI29.MM28_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI31.MM28 N_XI13.XI31.NET31_XI13.XI31.MM28_d
+ N_XI13.XI31.CLKB_XI13.XI31.MM28_g N_XI13.XI31.NET58_XI13.XI31.MM28_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI28.MM28 N_XI13.XI28.NET31_XI13.XI28.MM28_d
+ N_XI13.XI28.CLKB_XI13.XI28.MM28_g N_XI13.XI28.NET58_XI13.XI28.MM28_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI25.MM28 N_XI13.XI25.NET31_XI13.XI25.MM28_d
+ N_XI13.XI25.CLKB_XI13.XI25.MM28_g N_XI13.XI25.NET58_XI13.XI25.MM28_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI26.MM28 N_XI13.XI26.NET31_XI13.XI26.MM28_d
+ N_XI13.XI26.CLKB_XI13.XI26.MM28_g N_XI13.XI26.NET58_XI13.XI26.MM28_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI24.MM28 N_XI13.XI24.NET31_XI13.XI24.MM28_d
+ N_XI13.XI24.CLKB_XI13.XI24.MM28_g N_XI13.XI24.NET58_XI13.XI24.MM28_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI27.MM28 N_XI13.XI27.NET31_XI13.XI27.MM28_d
+ N_XI13.XI27.CLKB_XI13.XI27.MM28_g N_XI13.XI27.NET58_XI13.XI27.MM28_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI22.MM28 N_XI13.XI22.NET31_XI13.XI22.MM28_d
+ N_XI13.XI22.CLKB_XI13.XI22.MM28_g N_XI13.XI22.NET58_XI13.XI22.MM28_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI21.MM28 N_XI13.XI21.NET31_XI13.XI21.MM28_d
+ N_XI13.XI21.CLKB_XI13.XI21.MM28_g N_XI13.XI21.NET58_XI13.XI21.MM28_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI23.MM28 N_XI13.XI23.NET31_XI13.XI23.MM28_d
+ N_XI13.XI23.CLKB_XI13.XI23.MM28_g N_XI13.XI23.NET58_XI13.XI23.MM28_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI19.MM28 N_XI13.XI19.NET31_XI13.XI19.MM28_d
+ N_XI13.XI19.CLKB_XI13.XI19.MM28_g N_XI13.XI19.NET58_XI13.XI19.MM28_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI20.MM28 N_XI13.XI20.NET31_XI13.XI20.MM28_d
+ N_XI13.XI20.CLKB_XI13.XI20.MM28_g N_XI13.XI20.NET58_XI13.XI20.MM28_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI18.MM28 N_XI13.XI18.NET31_XI13.XI18.MM28_d
+ N_XI13.XI18.CLKB_XI13.XI18.MM28_g N_XI13.XI18.NET58_XI13.XI18.MM28_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI17.MM28 N_XI13.XI17.NET31_XI13.XI17.MM28_d
+ N_XI13.XI17.CLKB_XI13.XI17.MM28_g N_XI13.XI17.NET58_XI13.XI17.MM28_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI0.MM28 N_XI13.XI0.NET31_XI13.XI0.MM28_d N_XI13.XI0.CLKB_XI13.XI0.MM28_g
+ N_XI13.XI0.NET58_XI13.XI0.MM28_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI13.XI30.MM6 N_XI13.XI30.NET15_XI13.XI30.MM6_d
+ N_XI13.XI30.NET58_XI13.XI30.MM6_g N_VSS_XI13.XI30.MM6_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI29.MM6 N_XI13.XI29.NET15_XI13.XI29.MM6_d
+ N_XI13.XI29.NET58_XI13.XI29.MM6_g N_VSS_XI13.XI29.MM6_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI31.MM6 N_XI13.XI31.NET15_XI13.XI31.MM6_d
+ N_XI13.XI31.NET58_XI13.XI31.MM6_g N_VSS_XI13.XI31.MM6_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI28.MM6 N_XI13.XI28.NET15_XI13.XI28.MM6_d
+ N_XI13.XI28.NET58_XI13.XI28.MM6_g N_VSS_XI13.XI28.MM6_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI25.MM6 N_XI13.XI25.NET15_XI13.XI25.MM6_d
+ N_XI13.XI25.NET58_XI13.XI25.MM6_g N_VSS_XI13.XI25.MM6_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI26.MM6 N_XI13.XI26.NET15_XI13.XI26.MM6_d
+ N_XI13.XI26.NET58_XI13.XI26.MM6_g N_VSS_XI13.XI26.MM6_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI24.MM6 N_XI13.XI24.NET15_XI13.XI24.MM6_d
+ N_XI13.XI24.NET58_XI13.XI24.MM6_g N_VSS_XI13.XI24.MM6_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI27.MM6 N_XI13.XI27.NET15_XI13.XI27.MM6_d
+ N_XI13.XI27.NET58_XI13.XI27.MM6_g N_VSS_XI13.XI27.MM6_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI22.MM6 N_XI13.XI22.NET15_XI13.XI22.MM6_d
+ N_XI13.XI22.NET58_XI13.XI22.MM6_g N_VSS_XI13.XI22.MM6_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI21.MM6 N_XI13.XI21.NET15_XI13.XI21.MM6_d
+ N_XI13.XI21.NET58_XI13.XI21.MM6_g N_VSS_XI13.XI21.MM6_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI23.MM6 N_XI13.XI23.NET15_XI13.XI23.MM6_d
+ N_XI13.XI23.NET58_XI13.XI23.MM6_g N_VSS_XI13.XI23.MM6_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI19.MM6 N_XI13.XI19.NET15_XI13.XI19.MM6_d
+ N_XI13.XI19.NET58_XI13.XI19.MM6_g N_VSS_XI13.XI19.MM6_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI20.MM6 N_XI13.XI20.NET15_XI13.XI20.MM6_d
+ N_XI13.XI20.NET58_XI13.XI20.MM6_g N_VSS_XI13.XI20.MM6_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI18.MM6 N_XI13.XI18.NET15_XI13.XI18.MM6_d
+ N_XI13.XI18.NET58_XI13.XI18.MM6_g N_VSS_XI13.XI18.MM6_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI17.MM6 N_XI13.XI17.NET15_XI13.XI17.MM6_d
+ N_XI13.XI17.NET58_XI13.XI17.MM6_g N_VSS_XI13.XI17.MM6_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI0.MM6 N_XI13.XI0.NET15_XI13.XI0.MM6_d N_XI13.XI0.NET58_XI13.XI0.MM6_g
+ N_VSS_XI13.XI0.MM6_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI13.XI30.MM0 N_XI13.XI30.NET54_XI13.XI30.MM0_d
+ N_XI13.XI30.NET15_XI13.XI30.MM0_g N_VSS_XI13.XI30.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI29.MM0 N_XI13.XI29.NET54_XI13.XI29.MM0_d
+ N_XI13.XI29.NET15_XI13.XI29.MM0_g N_VSS_XI13.XI29.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI31.MM0 N_XI13.XI31.NET54_XI13.XI31.MM0_d
+ N_XI13.XI31.NET15_XI13.XI31.MM0_g N_VSS_XI13.XI31.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI28.MM0 N_XI13.XI28.NET54_XI13.XI28.MM0_d
+ N_XI13.XI28.NET15_XI13.XI28.MM0_g N_VSS_XI13.XI28.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI25.MM0 N_XI13.XI25.NET54_XI13.XI25.MM0_d
+ N_XI13.XI25.NET15_XI13.XI25.MM0_g N_VSS_XI13.XI25.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI26.MM0 N_XI13.XI26.NET54_XI13.XI26.MM0_d
+ N_XI13.XI26.NET15_XI13.XI26.MM0_g N_VSS_XI13.XI26.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI24.MM0 N_XI13.XI24.NET54_XI13.XI24.MM0_d
+ N_XI13.XI24.NET15_XI13.XI24.MM0_g N_VSS_XI13.XI24.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI27.MM0 N_XI13.XI27.NET54_XI13.XI27.MM0_d
+ N_XI13.XI27.NET15_XI13.XI27.MM0_g N_VSS_XI13.XI27.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI22.MM0 N_XI13.XI22.NET54_XI13.XI22.MM0_d
+ N_XI13.XI22.NET15_XI13.XI22.MM0_g N_VSS_XI13.XI22.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI21.MM0 N_XI13.XI21.NET54_XI13.XI21.MM0_d
+ N_XI13.XI21.NET15_XI13.XI21.MM0_g N_VSS_XI13.XI21.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI23.MM0 N_XI13.XI23.NET54_XI13.XI23.MM0_d
+ N_XI13.XI23.NET15_XI13.XI23.MM0_g N_VSS_XI13.XI23.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI19.MM0 N_XI13.XI19.NET54_XI13.XI19.MM0_d
+ N_XI13.XI19.NET15_XI13.XI19.MM0_g N_VSS_XI13.XI19.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI20.MM0 N_XI13.XI20.NET54_XI13.XI20.MM0_d
+ N_XI13.XI20.NET15_XI13.XI20.MM0_g N_VSS_XI13.XI20.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI18.MM0 N_XI13.XI18.NET54_XI13.XI18.MM0_d
+ N_XI13.XI18.NET15_XI13.XI18.MM0_g N_VSS_XI13.XI18.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI17.MM0 N_XI13.XI17.NET54_XI13.XI17.MM0_d
+ N_XI13.XI17.NET15_XI13.XI17.MM0_g N_VSS_XI13.XI17.MM0_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI0.MM0 N_XI13.XI0.NET54_XI13.XI0.MM0_d N_XI13.XI0.NET15_XI13.XI0.MM0_g
+ N_VSS_XI13.XI0.MM0_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI13.XI30.MM36 N_XI13.XI30.NET58_XI13.XI30.MM36_d
+ N_XI13.XI30.NET35_XI13.XI30.MM36_g N_XI13.XI30.NET54_XI13.XI30.MM36_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI29.MM36 N_XI13.XI29.NET58_XI13.XI29.MM36_d
+ N_XI13.XI29.NET35_XI13.XI29.MM36_g N_XI13.XI29.NET54_XI13.XI29.MM36_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI31.MM36 N_XI13.XI31.NET58_XI13.XI31.MM36_d
+ N_XI13.XI31.NET35_XI13.XI31.MM36_g N_XI13.XI31.NET54_XI13.XI31.MM36_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI28.MM36 N_XI13.XI28.NET58_XI13.XI28.MM36_d
+ N_XI13.XI28.NET35_XI13.XI28.MM36_g N_XI13.XI28.NET54_XI13.XI28.MM36_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI25.MM36 N_XI13.XI25.NET58_XI13.XI25.MM36_d
+ N_XI13.XI25.NET35_XI13.XI25.MM36_g N_XI13.XI25.NET54_XI13.XI25.MM36_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI26.MM36 N_XI13.XI26.NET58_XI13.XI26.MM36_d
+ N_XI13.XI26.NET35_XI13.XI26.MM36_g N_XI13.XI26.NET54_XI13.XI26.MM36_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI24.MM36 N_XI13.XI24.NET58_XI13.XI24.MM36_d
+ N_XI13.XI24.NET35_XI13.XI24.MM36_g N_XI13.XI24.NET54_XI13.XI24.MM36_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI27.MM36 N_XI13.XI27.NET58_XI13.XI27.MM36_d
+ N_XI13.XI27.NET35_XI13.XI27.MM36_g N_XI13.XI27.NET54_XI13.XI27.MM36_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI22.MM36 N_XI13.XI22.NET58_XI13.XI22.MM36_d
+ N_XI13.XI22.NET35_XI13.XI22.MM36_g N_XI13.XI22.NET54_XI13.XI22.MM36_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI21.MM36 N_XI13.XI21.NET58_XI13.XI21.MM36_d
+ N_XI13.XI21.NET35_XI13.XI21.MM36_g N_XI13.XI21.NET54_XI13.XI21.MM36_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI23.MM36 N_XI13.XI23.NET58_XI13.XI23.MM36_d
+ N_XI13.XI23.NET35_XI13.XI23.MM36_g N_XI13.XI23.NET54_XI13.XI23.MM36_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI19.MM36 N_XI13.XI19.NET58_XI13.XI19.MM36_d
+ N_XI13.XI19.NET35_XI13.XI19.MM36_g N_XI13.XI19.NET54_XI13.XI19.MM36_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI20.MM36 N_XI13.XI20.NET58_XI13.XI20.MM36_d
+ N_XI13.XI20.NET35_XI13.XI20.MM36_g N_XI13.XI20.NET54_XI13.XI20.MM36_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI18.MM36 N_XI13.XI18.NET58_XI13.XI18.MM36_d
+ N_XI13.XI18.NET35_XI13.XI18.MM36_g N_XI13.XI18.NET54_XI13.XI18.MM36_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI17.MM36 N_XI13.XI17.NET58_XI13.XI17.MM36_d
+ N_XI13.XI17.NET35_XI13.XI17.MM36_g N_XI13.XI17.NET54_XI13.XI17.MM36_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI0.MM36 N_XI13.XI0.NET58_XI13.XI0.MM36_d N_XI13.XI0.NET35_XI13.XI0.MM36_g
+ N_XI13.XI0.NET54_XI13.XI0.MM36_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI13.XI30.MM38 N_XI13.XI30.NET15_XI13.XI30.MM38_d
+ N_XI13.XI30.NET35_XI13.XI30.MM38_g N_XI13.XI30.NET14_XI13.XI30.MM38_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI29.MM38 N_XI13.XI29.NET15_XI13.XI29.MM38_d
+ N_XI13.XI29.NET35_XI13.XI29.MM38_g N_XI13.XI29.NET14_XI13.XI29.MM38_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI31.MM38 N_XI13.XI31.NET15_XI13.XI31.MM38_d
+ N_XI13.XI31.NET35_XI13.XI31.MM38_g N_XI13.XI31.NET14_XI13.XI31.MM38_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI28.MM38 N_XI13.XI28.NET15_XI13.XI28.MM38_d
+ N_XI13.XI28.NET35_XI13.XI28.MM38_g N_XI13.XI28.NET14_XI13.XI28.MM38_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI25.MM38 N_XI13.XI25.NET15_XI13.XI25.MM38_d
+ N_XI13.XI25.NET35_XI13.XI25.MM38_g N_XI13.XI25.NET14_XI13.XI25.MM38_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI26.MM38 N_XI13.XI26.NET15_XI13.XI26.MM38_d
+ N_XI13.XI26.NET35_XI13.XI26.MM38_g N_XI13.XI26.NET14_XI13.XI26.MM38_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI24.MM38 N_XI13.XI24.NET15_XI13.XI24.MM38_d
+ N_XI13.XI24.NET35_XI13.XI24.MM38_g N_XI13.XI24.NET14_XI13.XI24.MM38_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI27.MM38 N_XI13.XI27.NET15_XI13.XI27.MM38_d
+ N_XI13.XI27.NET35_XI13.XI27.MM38_g N_XI13.XI27.NET14_XI13.XI27.MM38_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI22.MM38 N_XI13.XI22.NET15_XI13.XI22.MM38_d
+ N_XI13.XI22.NET35_XI13.XI22.MM38_g N_XI13.XI22.NET14_XI13.XI22.MM38_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI21.MM38 N_XI13.XI21.NET15_XI13.XI21.MM38_d
+ N_XI13.XI21.NET35_XI13.XI21.MM38_g N_XI13.XI21.NET14_XI13.XI21.MM38_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI23.MM38 N_XI13.XI23.NET15_XI13.XI23.MM38_d
+ N_XI13.XI23.NET35_XI13.XI23.MM38_g N_XI13.XI23.NET14_XI13.XI23.MM38_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI19.MM38 N_XI13.XI19.NET15_XI13.XI19.MM38_d
+ N_XI13.XI19.NET35_XI13.XI19.MM38_g N_XI13.XI19.NET14_XI13.XI19.MM38_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI20.MM38 N_XI13.XI20.NET15_XI13.XI20.MM38_d
+ N_XI13.XI20.NET35_XI13.XI20.MM38_g N_XI13.XI20.NET14_XI13.XI20.MM38_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI18.MM38 N_XI13.XI18.NET15_XI13.XI18.MM38_d
+ N_XI13.XI18.NET35_XI13.XI18.MM38_g N_XI13.XI18.NET14_XI13.XI18.MM38_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI17.MM38 N_XI13.XI17.NET15_XI13.XI17.MM38_d
+ N_XI13.XI17.NET35_XI13.XI17.MM38_g N_XI13.XI17.NET14_XI13.XI17.MM38_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI0.MM38 N_XI13.XI0.NET15_XI13.XI0.MM38_d N_XI13.XI0.NET35_XI13.XI0.MM38_g
+ N_XI13.XI0.NET14_XI13.XI0.MM38_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI13.XI30.MM15 N_MAX15_XI13.XI30.MM15_d N_XI13.XI30.NET14_XI13.XI30.MM15_g
+ N_VSS_XI13.XI30.MM15_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI13.XI29.MM15 N_MAX14_XI13.XI29.MM15_d N_XI13.XI29.NET14_XI13.XI29.MM15_g
+ N_VSS_XI13.XI29.MM15_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI13.XI31.MM15 N_MAX13_XI13.XI31.MM15_d N_XI13.XI31.NET14_XI13.XI31.MM15_g
+ N_VSS_XI13.XI31.MM15_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI13.XI28.MM15 N_MAX12_XI13.XI28.MM15_d N_XI13.XI28.NET14_XI13.XI28.MM15_g
+ N_VSS_XI13.XI28.MM15_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI13.XI25.MM15 N_MAX11_XI13.XI25.MM15_d N_XI13.XI25.NET14_XI13.XI25.MM15_g
+ N_VSS_XI13.XI25.MM15_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI13.XI26.MM15 N_MAX10_XI13.XI26.MM15_d N_XI13.XI26.NET14_XI13.XI26.MM15_g
+ N_VSS_XI13.XI26.MM15_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI13.XI24.MM15 N_MAX9_XI13.XI24.MM15_d N_XI13.XI24.NET14_XI13.XI24.MM15_g
+ N_VSS_XI13.XI24.MM15_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI13.XI27.MM15 N_MAX8_XI13.XI27.MM15_d N_XI13.XI27.NET14_XI13.XI27.MM15_g
+ N_VSS_XI13.XI27.MM15_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI13.XI22.MM15 N_MAX7_XI13.XI22.MM15_d N_XI13.XI22.NET14_XI13.XI22.MM15_g
+ N_VSS_XI13.XI22.MM15_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI13.XI21.MM15 N_MAX6_XI13.XI21.MM15_d N_XI13.XI21.NET14_XI13.XI21.MM15_g
+ N_VSS_XI13.XI21.MM15_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI13.XI23.MM15 N_MAX5_XI13.XI23.MM15_d N_XI13.XI23.NET14_XI13.XI23.MM15_g
+ N_VSS_XI13.XI23.MM15_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI13.XI19.MM15 N_MAX4_XI13.XI19.MM15_d N_XI13.XI19.NET14_XI13.XI19.MM15_g
+ N_VSS_XI13.XI19.MM15_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI13.XI20.MM15 N_MAX3_XI13.XI20.MM15_d N_XI13.XI20.NET14_XI13.XI20.MM15_g
+ N_VSS_XI13.XI20.MM15_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI13.XI18.MM15 N_MAX2_XI13.XI18.MM15_d N_XI13.XI18.NET14_XI13.XI18.MM15_g
+ N_VSS_XI13.XI18.MM15_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI13.XI17.MM15 N_MAX1_XI13.XI17.MM15_d N_XI13.XI17.NET14_XI13.XI17.MM15_g
+ N_VSS_XI13.XI17.MM15_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI13.XI0.MM15 N_MAX0_XI13.XI0.MM15_d N_XI13.XI0.NET14_XI13.XI0.MM15_g
+ N_VSS_XI13.XI0.MM15_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI13.XI30.MM16 N_XI13.BAR_Q16_XI13.XI30.MM16_d N_MAX15_XI13.XI30.MM16_g
+ N_VSS_XI13.XI30.MM16_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI13.XI29.MM16 N_XI13.BAR_Q15_XI13.XI29.MM16_d N_MAX14_XI13.XI29.MM16_g
+ N_VSS_XI13.XI29.MM16_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI13.XI31.MM16 N_XI13.BAR_Q14_XI13.XI31.MM16_d N_MAX13_XI13.XI31.MM16_g
+ N_VSS_XI13.XI31.MM16_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI13.XI28.MM16 N_XI13.BAR_Q13_XI13.XI28.MM16_d N_MAX12_XI13.XI28.MM16_g
+ N_VSS_XI13.XI28.MM16_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI13.XI25.MM16 N_XI13.BAR_Q12_XI13.XI25.MM16_d N_MAX11_XI13.XI25.MM16_g
+ N_VSS_XI13.XI25.MM16_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI13.XI26.MM16 N_XI13.BAR_Q11_XI13.XI26.MM16_d N_MAX10_XI13.XI26.MM16_g
+ N_VSS_XI13.XI26.MM16_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI13.XI24.MM16 N_XI13.BAR_Q10_XI13.XI24.MM16_d N_MAX9_XI13.XI24.MM16_g
+ N_VSS_XI13.XI24.MM16_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI13.XI27.MM16 N_XI13.BAR_Q9_XI13.XI27.MM16_d N_MAX8_XI13.XI27.MM16_g
+ N_VSS_XI13.XI27.MM16_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI13.XI22.MM16 N_XI13.BAR_Q8_XI13.XI22.MM16_d N_MAX7_XI13.XI22.MM16_g
+ N_VSS_XI13.XI22.MM16_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI13.XI21.MM16 N_XI13.BAR_Q7_XI13.XI21.MM16_d N_MAX6_XI13.XI21.MM16_g
+ N_VSS_XI13.XI21.MM16_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI13.XI23.MM16 N_XI13.BAR_Q6_XI13.XI23.MM16_d N_MAX5_XI13.XI23.MM16_g
+ N_VSS_XI13.XI23.MM16_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI13.XI19.MM16 N_XI13.BAR_Q5_XI13.XI19.MM16_d N_MAX4_XI13.XI19.MM16_g
+ N_VSS_XI13.XI19.MM16_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI13.XI20.MM16 N_XI13.BAR_Q4_XI13.XI20.MM16_d N_MAX3_XI13.XI20.MM16_g
+ N_VSS_XI13.XI20.MM16_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI13.XI18.MM16 N_XI13.BAR_Q3_XI13.XI18.MM16_d N_MAX2_XI13.XI18.MM16_g
+ N_VSS_XI13.XI18.MM16_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI13.XI17.MM16 N_XI13.BAR_Q2_XI13.XI17.MM16_d N_MAX1_XI13.XI17.MM16_g
+ N_VSS_XI13.XI17.MM16_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI13.XI0.MM16 N_XI13.BAR_Q1_XI13.XI0.MM16_d N_MAX0_XI13.XI0.MM16_g
+ N_VSS_XI13.XI0.MM16_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI13.XI30.MM40 N_XI13.XI30.NET14_XI13.XI30.MM40_d
+ N_XI13.XI30.CLKB_XI13.XI30.MM40_g N_XI13.BAR_Q16_XI13.XI30.MM40_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI29.MM40 N_XI13.XI29.NET14_XI13.XI29.MM40_d
+ N_XI13.XI29.CLKB_XI13.XI29.MM40_g N_XI13.BAR_Q15_XI13.XI29.MM40_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI31.MM40 N_XI13.XI31.NET14_XI13.XI31.MM40_d
+ N_XI13.XI31.CLKB_XI13.XI31.MM40_g N_XI13.BAR_Q14_XI13.XI31.MM40_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI28.MM40 N_XI13.XI28.NET14_XI13.XI28.MM40_d
+ N_XI13.XI28.CLKB_XI13.XI28.MM40_g N_XI13.BAR_Q13_XI13.XI28.MM40_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI25.MM40 N_XI13.XI25.NET14_XI13.XI25.MM40_d
+ N_XI13.XI25.CLKB_XI13.XI25.MM40_g N_XI13.BAR_Q12_XI13.XI25.MM40_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI26.MM40 N_XI13.XI26.NET14_XI13.XI26.MM40_d
+ N_XI13.XI26.CLKB_XI13.XI26.MM40_g N_XI13.BAR_Q11_XI13.XI26.MM40_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI24.MM40 N_XI13.XI24.NET14_XI13.XI24.MM40_d
+ N_XI13.XI24.CLKB_XI13.XI24.MM40_g N_XI13.BAR_Q10_XI13.XI24.MM40_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI27.MM40 N_XI13.XI27.NET14_XI13.XI27.MM40_d
+ N_XI13.XI27.CLKB_XI13.XI27.MM40_g N_XI13.BAR_Q9_XI13.XI27.MM40_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI22.MM40 N_XI13.XI22.NET14_XI13.XI22.MM40_d
+ N_XI13.XI22.CLKB_XI13.XI22.MM40_g N_XI13.BAR_Q8_XI13.XI22.MM40_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI21.MM40 N_XI13.XI21.NET14_XI13.XI21.MM40_d
+ N_XI13.XI21.CLKB_XI13.XI21.MM40_g N_XI13.BAR_Q7_XI13.XI21.MM40_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI23.MM40 N_XI13.XI23.NET14_XI13.XI23.MM40_d
+ N_XI13.XI23.CLKB_XI13.XI23.MM40_g N_XI13.BAR_Q6_XI13.XI23.MM40_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI19.MM40 N_XI13.XI19.NET14_XI13.XI19.MM40_d
+ N_XI13.XI19.CLKB_XI13.XI19.MM40_g N_XI13.BAR_Q5_XI13.XI19.MM40_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI20.MM40 N_XI13.XI20.NET14_XI13.XI20.MM40_d
+ N_XI13.XI20.CLKB_XI13.XI20.MM40_g N_XI13.BAR_Q4_XI13.XI20.MM40_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI18.MM40 N_XI13.XI18.NET14_XI13.XI18.MM40_d
+ N_XI13.XI18.CLKB_XI13.XI18.MM40_g N_XI13.BAR_Q3_XI13.XI18.MM40_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI17.MM40 N_XI13.XI17.NET14_XI13.XI17.MM40_d
+ N_XI13.XI17.CLKB_XI13.XI17.MM40_g N_XI13.BAR_Q2_XI13.XI17.MM40_s
+ N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07 AD=3.75e-13 AS=3.75e-13
+ PD=2e-06 PS=2e-06
mXI13.XI0.MM40 N_XI13.XI0.NET14_XI13.XI0.MM40_d N_XI13.XI0.CLKB_XI13.XI0.MM40_g
+ N_XI13.BAR_Q1_XI13.XI0.MM40_s N_VSS_XI10.XI0.XI0.MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=3.75e-13 AS=3.75e-13 PD=2e-06 PS=2e-06
mXI10.XI0.XI0.MM1 N_XI10.XI0.NET0180_XI10.XI0.XI0.MM1_d
+ N_NET222_XI10.XI0.XI0.MM1_g N_VDD_XI10.XI0.XI0.MM1_s N_VDD_XI10.XI0.XI0.MM1_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI25.MM1 N_NET206_XI25.MM1_d N_CLEAR_XI25.MM1_g N_VDD_XI25.MM1_s
+ N_VDD_XI25.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06
+ PS=2.48e-06
mXI24.MM1 N_NET202_XI24.MM1_d N_NET206_XI24.MM1_g N_VDD_XI24.MM1_s
+ N_VDD_XI25.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06
+ PS=2.48e-06
mXI23.XI11.MM1 N_NET696_XI23.XI11.MM1_d N_A15_XI23.XI11.MM1_g
+ N_VDD_XI23.XI11.MM1_s N_VDD_XI23.XI11.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI22.XI11.MM1 N_NET662_XI22.XI11.MM1_d N_NET696_XI22.XI11.MM1_g
+ N_VDD_XI22.XI11.MM1_s N_VDD_XI23.XI11.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI23.XI12.MM1 N_NET697_XI23.XI12.MM1_d N_A14_XI23.XI12.MM1_g
+ N_VDD_XI23.XI12.MM1_s N_VDD_XI23.XI11.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI22.XI12.MM1 N_NET663_XI22.XI12.MM1_d N_NET697_XI22.XI12.MM1_g
+ N_VDD_XI22.XI12.MM1_s N_VDD_XI23.XI11.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI23.XI10.MM1 N_NET698_XI23.XI10.MM1_d N_A13_XI23.XI10.MM1_g
+ N_VDD_XI23.XI10.MM1_s N_VDD_XI23.XI11.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI22.XI10.MM1 N_NET664_XI22.XI10.MM1_d N_NET698_XI22.XI10.MM1_g
+ N_VDD_XI22.XI10.MM1_s N_VDD_XI23.XI11.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI23.XI9.MM1 N_NET699_XI23.XI9.MM1_d N_A12_XI23.XI9.MM1_g N_VDD_XI23.XI9.MM1_s
+ N_VDD_XI23.XI11.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI22.XI9.MM1 N_NET665_XI22.XI9.MM1_d N_NET699_XI22.XI9.MM1_g
+ N_VDD_XI22.XI9.MM1_s N_VDD_XI23.XI11.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI23.XI14.MM1 N_NET700_XI23.XI14.MM1_d N_A11_XI23.XI14.MM1_g
+ N_VDD_XI23.XI14.MM1_s N_VDD_XI23.XI11.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI22.XI14.MM1 N_NET666_XI22.XI14.MM1_d N_NET700_XI22.XI14.MM1_g
+ N_VDD_XI22.XI14.MM1_s N_VDD_XI23.XI11.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI23.XI13.MM1 N_NET701_XI23.XI13.MM1_d N_A10_XI23.XI13.MM1_g
+ N_VDD_XI23.XI13.MM1_s N_VDD_XI23.XI11.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI22.XI13.MM1 N_NET667_XI22.XI13.MM1_d N_NET701_XI22.XI13.MM1_g
+ N_VDD_XI22.XI13.MM1_s N_VDD_XI23.XI11.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI23.XI15.MM1 N_NET702_XI23.XI15.MM1_d N_A9_XI23.XI15.MM1_g
+ N_VDD_XI23.XI15.MM1_s N_VDD_XI23.XI11.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI22.XI15.MM1 N_NET668_XI22.XI15.MM1_d N_NET702_XI22.XI15.MM1_g
+ N_VDD_XI22.XI15.MM1_s N_VDD_XI23.XI11.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI23.XI6.MM1 N_NET703_XI23.XI6.MM1_d N_A8_XI23.XI6.MM1_g N_VDD_XI23.XI6.MM1_s
+ N_VDD_XI23.XI11.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI22.XI6.MM1 N_NET669_XI22.XI6.MM1_d N_NET703_XI22.XI6.MM1_g
+ N_VDD_XI22.XI6.MM1_s N_VDD_XI23.XI11.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI23.XI5.MM1 N_NET704_XI23.XI5.MM1_d N_A7_XI23.XI5.MM1_g N_VDD_XI23.XI5.MM1_s
+ N_VDD_XI23.XI11.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI22.XI5.MM1 N_NET670_XI22.XI5.MM1_d N_NET704_XI22.XI5.MM1_g
+ N_VDD_XI22.XI5.MM1_s N_VDD_XI23.XI11.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI23.XI7.MM1 N_NET705_XI23.XI7.MM1_d N_A6_XI23.XI7.MM1_g N_VDD_XI23.XI7.MM1_s
+ N_VDD_XI23.XI11.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI22.XI7.MM1 N_NET671_XI22.XI7.MM1_d N_NET705_XI22.XI7.MM1_g
+ N_VDD_XI22.XI7.MM1_s N_VDD_XI23.XI11.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI23.XI8.MM1 N_NET706_XI23.XI8.MM1_d N_A5_XI23.XI8.MM1_g N_VDD_XI23.XI8.MM1_s
+ N_VDD_XI23.XI11.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI22.XI8.MM1 N_NET672_XI22.XI8.MM1_d N_NET706_XI22.XI8.MM1_g
+ N_VDD_XI22.XI8.MM1_s N_VDD_XI23.XI11.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI23.XI3.MM1 N_NET707_XI23.XI3.MM1_d N_A4_XI23.XI3.MM1_g N_VDD_XI23.XI3.MM1_s
+ N_VDD_XI23.XI11.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI22.XI3.MM1 N_NET673_XI22.XI3.MM1_d N_NET707_XI22.XI3.MM1_g
+ N_VDD_XI22.XI3.MM1_s N_VDD_XI23.XI11.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI23.XI4.MM1 N_NET708_XI23.XI4.MM1_d N_A3_XI23.XI4.MM1_g N_VDD_XI23.XI4.MM1_s
+ N_VDD_XI23.XI11.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI22.XI4.MM1 N_NET674_XI22.XI4.MM1_d N_NET708_XI22.XI4.MM1_g
+ N_VDD_XI22.XI4.MM1_s N_VDD_XI23.XI11.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI23.XI2.MM1 N_NET709_XI23.XI2.MM1_d N_A2_XI23.XI2.MM1_g N_VDD_XI23.XI2.MM1_s
+ N_VDD_XI23.XI11.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI22.XI2.MM1 N_NET675_XI22.XI2.MM1_d N_NET709_XI22.XI2.MM1_g
+ N_VDD_XI22.XI2.MM1_s N_VDD_XI23.XI11.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI23.XI1.MM1 N_NET710_XI23.XI1.MM1_d N_A1_XI23.XI1.MM1_g N_VDD_XI23.XI1.MM1_s
+ N_VDD_XI23.XI11.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI22.XI1.MM1 N_NET676_XI22.XI1.MM1_d N_NET710_XI22.XI1.MM1_g
+ N_VDD_XI22.XI1.MM1_s N_VDD_XI23.XI11.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI23.XI0.MM1 N_NET711_XI23.XI0.MM1_d N_A0_XI23.XI0.MM1_g N_VDD_XI23.XI0.MM1_s
+ N_VDD_XI23.XI11.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI22.XI0.MM1 N_NET677_XI22.XI0.MM1_d N_NET711_XI22.XI0.MM1_g
+ N_VDD_XI22.XI0.MM1_s N_VDD_XI23.XI11.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI17.MM35 N_XI17.NET58_XI17.MM35_d N_XI17.CLKB_XI17.MM35_g
+ N_XI17.NET54_XI17.MM35_s N_VDD_XI17.MM35_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI17.MM37 N_XI17.NET15_XI17.MM37_d N_XI17.CLKB_XI17.MM37_g
+ N_XI17.NET14_XI17.MM37_s N_VDD_XI17.MM35_b P_18 L=1.8e-07 W=1.5e-06
+ AD=1.125e-12 AS=9.375e-13 PD=3e-06 PS=2.75e-06
mXI17.MM39 N_XI17.NET14_XI17.MM39_d N_XI17.NET35_XI17.MM39_g
+ N_NET198_XI17.MM39_s N_VDD_XI17.MM35_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13
+ AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI17.XI0.MM1 N_XI17.NET0180_XI17.XI0.MM1_d N_NET222_XI17.XI0.MM1_g
+ N_VDD_XI17.XI0.MM1_s N_VDD_XI17.MM35_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13
+ AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI17.XI1.MM1 N_XI17.NET35_XI17.XI1.MM1_d N_XI17.NET0180_XI17.XI1.MM1_g
+ N_VDD_XI17.XI1.MM1_s N_VDD_XI17.MM35_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13
+ AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI17.MM25 N_XI17.CLKB_XI17.MM25_d N_XI17.NET35_XI17.MM25_g N_VDD_XI17.MM25_s
+ N_VDD_XI17.MM35_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI17.MM20 N_XI17.NET27_XI17.MM20_d N_NET202_XI17.MM20_g N_VDD_XI17.MM20_s
+ N_VDD_XI17.MM35_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI17.MM17 N_XI17.NET31_XI17.MM17_d N_XI17.NET27_XI17.MM17_g N_VDD_XI17.MM17_s
+ N_VDD_XI17.MM35_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI17.MM27 N_XI17.NET31_XI17.MM27_d N_XI17.NET35_XI17.MM27_g
+ N_XI17.NET58_XI17.MM27_s N_VDD_XI17.MM35_b P_18 L=1.8e-07 W=1.5e-06
+ AD=1.125e-12 AS=9.375e-13 PD=3e-06 PS=2.75e-06
mXI17.MM3 N_XI17.NET15_XI17.MM3_d N_XI17.NET58_XI17.MM3_g N_VDD_XI17.MM3_s
+ N_VDD_XI17.MM35_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI17.MM1 N_XI17.NET54_XI17.MM1_d N_XI17.NET15_XI17.MM1_g N_VDD_XI17.MM1_s
+ N_VDD_XI17.MM35_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI17.MM13 N_Q_XI17.MM13_d N_XI17.NET14_XI17.MM13_g N_VDD_XI17.MM13_s
+ N_VDD_XI17.MM35_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI17.MM14 N_NET198_XI17.MM14_d N_Q_XI17.MM14_g N_VDD_XI17.MM14_s
+ N_VDD_XI17.MM35_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI10.XI0.XI1.MM1 N_XI10.XI0.NET35_XI10.XI0.XI1.MM1_d
+ N_XI10.XI0.NET0180_XI10.XI0.XI1.MM1_g N_VDD_XI10.XI0.XI1.MM1_s
+ N_VDD_XI10.XI0.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI10.XI0.MM25 N_XI10.XI0.CLKB_XI10.XI0.MM25_d N_XI10.XI0.NET35_XI10.XI0.MM25_g
+ N_VDD_XI10.XI0.MM25_s N_VDD_XI10.XI0.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI10.XI0.MM20 N_XI10.XI0.NET27_XI10.XI0.MM20_d N_NET677_XI10.XI0.MM20_g
+ N_VDD_XI10.XI0.MM20_s N_VDD_XI10.XI0.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI10.XI0.MM17 N_XI10.XI0.NET31_XI10.XI0.MM17_d N_XI10.XI0.NET27_XI10.XI0.MM17_g
+ N_VDD_XI10.XI0.MM17_s N_VDD_XI10.XI0.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI10.XI30.XI0.MM1 N_XI10.XI30.NET0180_XI10.XI30.XI0.MM1_d
+ N_NET222_XI10.XI30.XI0.MM1_g N_VDD_XI10.XI30.XI0.MM1_s
+ N_VDD_XI10.XI30.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI10.XI29.XI0.MM1 N_XI10.XI29.NET0180_XI10.XI29.XI0.MM1_d
+ N_NET222_XI10.XI29.XI0.MM1_g N_VDD_XI10.XI29.XI0.MM1_s
+ N_VDD_XI10.XI29.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI10.XI31.XI0.MM1 N_XI10.XI31.NET0180_XI10.XI31.XI0.MM1_d
+ N_NET222_XI10.XI31.XI0.MM1_g N_VDD_XI10.XI31.XI0.MM1_s
+ N_VDD_XI10.XI31.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI10.XI28.XI0.MM1 N_XI10.XI28.NET0180_XI10.XI28.XI0.MM1_d
+ N_NET222_XI10.XI28.XI0.MM1_g N_VDD_XI10.XI28.XI0.MM1_s
+ N_VDD_XI10.XI28.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI10.XI25.XI0.MM1 N_XI10.XI25.NET0180_XI10.XI25.XI0.MM1_d
+ N_NET222_XI10.XI25.XI0.MM1_g N_VDD_XI10.XI25.XI0.MM1_s
+ N_VDD_XI10.XI25.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI10.XI26.XI0.MM1 N_XI10.XI26.NET0180_XI10.XI26.XI0.MM1_d
+ N_NET222_XI10.XI26.XI0.MM1_g N_VDD_XI10.XI26.XI0.MM1_s
+ N_VDD_XI10.XI26.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI10.XI24.XI0.MM1 N_XI10.XI24.NET0180_XI10.XI24.XI0.MM1_d
+ N_NET222_XI10.XI24.XI0.MM1_g N_VDD_XI10.XI24.XI0.MM1_s
+ N_VDD_XI10.XI24.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI10.XI27.XI0.MM1 N_XI10.XI27.NET0180_XI10.XI27.XI0.MM1_d
+ N_NET222_XI10.XI27.XI0.MM1_g N_VDD_XI10.XI27.XI0.MM1_s
+ N_VDD_XI10.XI27.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI10.XI22.XI0.MM1 N_XI10.XI22.NET0180_XI10.XI22.XI0.MM1_d
+ N_NET222_XI10.XI22.XI0.MM1_g N_VDD_XI10.XI22.XI0.MM1_s
+ N_VDD_XI10.XI22.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI10.XI21.XI0.MM1 N_XI10.XI21.NET0180_XI10.XI21.XI0.MM1_d
+ N_NET222_XI10.XI21.XI0.MM1_g N_VDD_XI10.XI21.XI0.MM1_s
+ N_VDD_XI10.XI21.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI10.XI23.XI0.MM1 N_XI10.XI23.NET0180_XI10.XI23.XI0.MM1_d
+ N_NET222_XI10.XI23.XI0.MM1_g N_VDD_XI10.XI23.XI0.MM1_s
+ N_VDD_XI10.XI23.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI10.XI19.XI0.MM1 N_XI10.XI19.NET0180_XI10.XI19.XI0.MM1_d
+ N_NET222_XI10.XI19.XI0.MM1_g N_VDD_XI10.XI19.XI0.MM1_s
+ N_VDD_XI10.XI19.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI10.XI20.XI0.MM1 N_XI10.XI20.NET0180_XI10.XI20.XI0.MM1_d
+ N_NET222_XI10.XI20.XI0.MM1_g N_VDD_XI10.XI20.XI0.MM1_s
+ N_VDD_XI10.XI20.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI10.XI18.XI0.MM1 N_XI10.XI18.NET0180_XI10.XI18.XI0.MM1_d
+ N_NET222_XI10.XI18.XI0.MM1_g N_VDD_XI10.XI18.XI0.MM1_s
+ N_VDD_XI10.XI18.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI10.XI17.XI0.MM1 N_XI10.XI17.NET0180_XI10.XI17.XI0.MM1_d
+ N_NET222_XI10.XI17.XI0.MM1_g N_VDD_XI10.XI17.XI0.MM1_s
+ N_VDD_XI10.XI17.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI10.XI0.MM27 N_XI10.XI0.NET31_XI10.XI0.MM27_d N_XI10.XI0.NET35_XI10.XI0.MM27_g
+ N_XI10.XI0.NET58_XI10.XI0.MM27_s N_VDD_XI10.XI0.XI0.MM1_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.125e-12 AS=9.375e-13 PD=3e-06 PS=2.75e-06
mXI10.XI30.XI1.MM1 N_XI10.XI30.NET35_XI10.XI30.XI1.MM1_d
+ N_XI10.XI30.NET0180_XI10.XI30.XI1.MM1_g N_VDD_XI10.XI30.XI1.MM1_s
+ N_VDD_XI10.XI30.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI10.XI29.XI1.MM1 N_XI10.XI29.NET35_XI10.XI29.XI1.MM1_d
+ N_XI10.XI29.NET0180_XI10.XI29.XI1.MM1_g N_VDD_XI10.XI29.XI1.MM1_s
+ N_VDD_XI10.XI29.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI10.XI31.XI1.MM1 N_XI10.XI31.NET35_XI10.XI31.XI1.MM1_d
+ N_XI10.XI31.NET0180_XI10.XI31.XI1.MM1_g N_VDD_XI10.XI31.XI1.MM1_s
+ N_VDD_XI10.XI31.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI10.XI28.XI1.MM1 N_XI10.XI28.NET35_XI10.XI28.XI1.MM1_d
+ N_XI10.XI28.NET0180_XI10.XI28.XI1.MM1_g N_VDD_XI10.XI28.XI1.MM1_s
+ N_VDD_XI10.XI28.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI10.XI25.XI1.MM1 N_XI10.XI25.NET35_XI10.XI25.XI1.MM1_d
+ N_XI10.XI25.NET0180_XI10.XI25.XI1.MM1_g N_VDD_XI10.XI25.XI1.MM1_s
+ N_VDD_XI10.XI25.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI10.XI26.XI1.MM1 N_XI10.XI26.NET35_XI10.XI26.XI1.MM1_d
+ N_XI10.XI26.NET0180_XI10.XI26.XI1.MM1_g N_VDD_XI10.XI26.XI1.MM1_s
+ N_VDD_XI10.XI26.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI10.XI24.XI1.MM1 N_XI10.XI24.NET35_XI10.XI24.XI1.MM1_d
+ N_XI10.XI24.NET0180_XI10.XI24.XI1.MM1_g N_VDD_XI10.XI24.XI1.MM1_s
+ N_VDD_XI10.XI24.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI10.XI27.XI1.MM1 N_XI10.XI27.NET35_XI10.XI27.XI1.MM1_d
+ N_XI10.XI27.NET0180_XI10.XI27.XI1.MM1_g N_VDD_XI10.XI27.XI1.MM1_s
+ N_VDD_XI10.XI27.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI10.XI22.XI1.MM1 N_XI10.XI22.NET35_XI10.XI22.XI1.MM1_d
+ N_XI10.XI22.NET0180_XI10.XI22.XI1.MM1_g N_VDD_XI10.XI22.XI1.MM1_s
+ N_VDD_XI10.XI22.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI10.XI21.XI1.MM1 N_XI10.XI21.NET35_XI10.XI21.XI1.MM1_d
+ N_XI10.XI21.NET0180_XI10.XI21.XI1.MM1_g N_VDD_XI10.XI21.XI1.MM1_s
+ N_VDD_XI10.XI21.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI10.XI23.XI1.MM1 N_XI10.XI23.NET35_XI10.XI23.XI1.MM1_d
+ N_XI10.XI23.NET0180_XI10.XI23.XI1.MM1_g N_VDD_XI10.XI23.XI1.MM1_s
+ N_VDD_XI10.XI23.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI10.XI19.XI1.MM1 N_XI10.XI19.NET35_XI10.XI19.XI1.MM1_d
+ N_XI10.XI19.NET0180_XI10.XI19.XI1.MM1_g N_VDD_XI10.XI19.XI1.MM1_s
+ N_VDD_XI10.XI19.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI10.XI20.XI1.MM1 N_XI10.XI20.NET35_XI10.XI20.XI1.MM1_d
+ N_XI10.XI20.NET0180_XI10.XI20.XI1.MM1_g N_VDD_XI10.XI20.XI1.MM1_s
+ N_VDD_XI10.XI20.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI10.XI18.XI1.MM1 N_XI10.XI18.NET35_XI10.XI18.XI1.MM1_d
+ N_XI10.XI18.NET0180_XI10.XI18.XI1.MM1_g N_VDD_XI10.XI18.XI1.MM1_s
+ N_VDD_XI10.XI18.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI10.XI17.XI1.MM1 N_XI10.XI17.NET35_XI10.XI17.XI1.MM1_d
+ N_XI10.XI17.NET0180_XI10.XI17.XI1.MM1_g N_VDD_XI10.XI17.XI1.MM1_s
+ N_VDD_XI10.XI17.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI10.XI0.MM3 N_XI10.XI0.NET15_XI10.XI0.MM3_d N_XI10.XI0.NET58_XI10.XI0.MM3_g
+ N_VDD_XI10.XI0.MM3_s N_VDD_XI10.XI0.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI10.XI30.MM25 N_XI10.XI30.CLKB_XI10.XI30.MM25_d
+ N_XI10.XI30.NET35_XI10.XI30.MM25_g N_VDD_XI10.XI30.MM25_s
+ N_VDD_XI10.XI30.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI10.XI29.MM25 N_XI10.XI29.CLKB_XI10.XI29.MM25_d
+ N_XI10.XI29.NET35_XI10.XI29.MM25_g N_VDD_XI10.XI29.MM25_s
+ N_VDD_XI10.XI29.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI10.XI31.MM25 N_XI10.XI31.CLKB_XI10.XI31.MM25_d
+ N_XI10.XI31.NET35_XI10.XI31.MM25_g N_VDD_XI10.XI31.MM25_s
+ N_VDD_XI10.XI31.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI10.XI28.MM25 N_XI10.XI28.CLKB_XI10.XI28.MM25_d
+ N_XI10.XI28.NET35_XI10.XI28.MM25_g N_VDD_XI10.XI28.MM25_s
+ N_VDD_XI10.XI28.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI10.XI25.MM25 N_XI10.XI25.CLKB_XI10.XI25.MM25_d
+ N_XI10.XI25.NET35_XI10.XI25.MM25_g N_VDD_XI10.XI25.MM25_s
+ N_VDD_XI10.XI25.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI10.XI26.MM25 N_XI10.XI26.CLKB_XI10.XI26.MM25_d
+ N_XI10.XI26.NET35_XI10.XI26.MM25_g N_VDD_XI10.XI26.MM25_s
+ N_VDD_XI10.XI26.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI10.XI24.MM25 N_XI10.XI24.CLKB_XI10.XI24.MM25_d
+ N_XI10.XI24.NET35_XI10.XI24.MM25_g N_VDD_XI10.XI24.MM25_s
+ N_VDD_XI10.XI24.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI10.XI27.MM25 N_XI10.XI27.CLKB_XI10.XI27.MM25_d
+ N_XI10.XI27.NET35_XI10.XI27.MM25_g N_VDD_XI10.XI27.MM25_s
+ N_VDD_XI10.XI27.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI10.XI22.MM25 N_XI10.XI22.CLKB_XI10.XI22.MM25_d
+ N_XI10.XI22.NET35_XI10.XI22.MM25_g N_VDD_XI10.XI22.MM25_s
+ N_VDD_XI10.XI22.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI10.XI21.MM25 N_XI10.XI21.CLKB_XI10.XI21.MM25_d
+ N_XI10.XI21.NET35_XI10.XI21.MM25_g N_VDD_XI10.XI21.MM25_s
+ N_VDD_XI10.XI21.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI10.XI23.MM25 N_XI10.XI23.CLKB_XI10.XI23.MM25_d
+ N_XI10.XI23.NET35_XI10.XI23.MM25_g N_VDD_XI10.XI23.MM25_s
+ N_VDD_XI10.XI23.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI10.XI19.MM25 N_XI10.XI19.CLKB_XI10.XI19.MM25_d
+ N_XI10.XI19.NET35_XI10.XI19.MM25_g N_VDD_XI10.XI19.MM25_s
+ N_VDD_XI10.XI19.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI10.XI20.MM25 N_XI10.XI20.CLKB_XI10.XI20.MM25_d
+ N_XI10.XI20.NET35_XI10.XI20.MM25_g N_VDD_XI10.XI20.MM25_s
+ N_VDD_XI10.XI20.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI10.XI18.MM25 N_XI10.XI18.CLKB_XI10.XI18.MM25_d
+ N_XI10.XI18.NET35_XI10.XI18.MM25_g N_VDD_XI10.XI18.MM25_s
+ N_VDD_XI10.XI18.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI10.XI17.MM25 N_XI10.XI17.CLKB_XI10.XI17.MM25_d
+ N_XI10.XI17.NET35_XI10.XI17.MM25_g N_VDD_XI10.XI17.MM25_s
+ N_VDD_XI10.XI17.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI10.XI0.MM1 N_XI10.XI0.NET54_XI10.XI0.MM1_d N_XI10.XI0.NET15_XI10.XI0.MM1_g
+ N_VDD_XI10.XI0.MM1_s N_VDD_XI10.XI0.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI10.XI30.MM20 N_XI10.XI30.NET27_XI10.XI30.MM20_d N_NET662_XI10.XI30.MM20_g
+ N_VDD_XI10.XI30.MM20_s N_VDD_XI10.XI30.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI10.XI29.MM20 N_XI10.XI29.NET27_XI10.XI29.MM20_d N_NET663_XI10.XI29.MM20_g
+ N_VDD_XI10.XI29.MM20_s N_VDD_XI10.XI29.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI10.XI31.MM20 N_XI10.XI31.NET27_XI10.XI31.MM20_d N_NET664_XI10.XI31.MM20_g
+ N_VDD_XI10.XI31.MM20_s N_VDD_XI10.XI31.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI10.XI28.MM20 N_XI10.XI28.NET27_XI10.XI28.MM20_d N_NET665_XI10.XI28.MM20_g
+ N_VDD_XI10.XI28.MM20_s N_VDD_XI10.XI28.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI10.XI25.MM20 N_XI10.XI25.NET27_XI10.XI25.MM20_d N_NET666_XI10.XI25.MM20_g
+ N_VDD_XI10.XI25.MM20_s N_VDD_XI10.XI25.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI10.XI26.MM20 N_XI10.XI26.NET27_XI10.XI26.MM20_d N_NET667_XI10.XI26.MM20_g
+ N_VDD_XI10.XI26.MM20_s N_VDD_XI10.XI26.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI10.XI24.MM20 N_XI10.XI24.NET27_XI10.XI24.MM20_d N_NET668_XI10.XI24.MM20_g
+ N_VDD_XI10.XI24.MM20_s N_VDD_XI10.XI24.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI10.XI27.MM20 N_XI10.XI27.NET27_XI10.XI27.MM20_d N_NET669_XI10.XI27.MM20_g
+ N_VDD_XI10.XI27.MM20_s N_VDD_XI10.XI27.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI10.XI22.MM20 N_XI10.XI22.NET27_XI10.XI22.MM20_d N_NET670_XI10.XI22.MM20_g
+ N_VDD_XI10.XI22.MM20_s N_VDD_XI10.XI22.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI10.XI21.MM20 N_XI10.XI21.NET27_XI10.XI21.MM20_d N_NET671_XI10.XI21.MM20_g
+ N_VDD_XI10.XI21.MM20_s N_VDD_XI10.XI21.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI10.XI23.MM20 N_XI10.XI23.NET27_XI10.XI23.MM20_d N_NET672_XI10.XI23.MM20_g
+ N_VDD_XI10.XI23.MM20_s N_VDD_XI10.XI23.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI10.XI19.MM20 N_XI10.XI19.NET27_XI10.XI19.MM20_d N_NET673_XI10.XI19.MM20_g
+ N_VDD_XI10.XI19.MM20_s N_VDD_XI10.XI19.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI10.XI20.MM20 N_XI10.XI20.NET27_XI10.XI20.MM20_d N_NET674_XI10.XI20.MM20_g
+ N_VDD_XI10.XI20.MM20_s N_VDD_XI10.XI20.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI10.XI18.MM20 N_XI10.XI18.NET27_XI10.XI18.MM20_d N_NET675_XI10.XI18.MM20_g
+ N_VDD_XI10.XI18.MM20_s N_VDD_XI10.XI18.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI10.XI17.MM20 N_XI10.XI17.NET27_XI10.XI17.MM20_d N_NET676_XI10.XI17.MM20_g
+ N_VDD_XI10.XI17.MM20_s N_VDD_XI10.XI17.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI10.XI0.MM35 N_XI10.XI0.NET58_XI10.XI0.MM35_d N_XI10.XI0.CLKB_XI10.XI0.MM35_g
+ N_XI10.XI0.NET54_XI10.XI0.MM35_s N_VDD_XI10.XI0.XI0.MM1_b P_18 L=1.8e-07
+ W=1.5e-06 AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI10.XI30.MM17 N_XI10.XI30.NET31_XI10.XI30.MM17_d
+ N_XI10.XI30.NET27_XI10.XI30.MM17_g N_VDD_XI10.XI30.MM17_s
+ N_VDD_XI10.XI30.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI10.XI29.MM17 N_XI10.XI29.NET31_XI10.XI29.MM17_d
+ N_XI10.XI29.NET27_XI10.XI29.MM17_g N_VDD_XI10.XI29.MM17_s
+ N_VDD_XI10.XI29.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI10.XI31.MM17 N_XI10.XI31.NET31_XI10.XI31.MM17_d
+ N_XI10.XI31.NET27_XI10.XI31.MM17_g N_VDD_XI10.XI31.MM17_s
+ N_VDD_XI10.XI31.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI10.XI28.MM17 N_XI10.XI28.NET31_XI10.XI28.MM17_d
+ N_XI10.XI28.NET27_XI10.XI28.MM17_g N_VDD_XI10.XI28.MM17_s
+ N_VDD_XI10.XI28.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI10.XI25.MM17 N_XI10.XI25.NET31_XI10.XI25.MM17_d
+ N_XI10.XI25.NET27_XI10.XI25.MM17_g N_VDD_XI10.XI25.MM17_s
+ N_VDD_XI10.XI25.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI10.XI26.MM17 N_XI10.XI26.NET31_XI10.XI26.MM17_d
+ N_XI10.XI26.NET27_XI10.XI26.MM17_g N_VDD_XI10.XI26.MM17_s
+ N_VDD_XI10.XI26.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI10.XI24.MM17 N_XI10.XI24.NET31_XI10.XI24.MM17_d
+ N_XI10.XI24.NET27_XI10.XI24.MM17_g N_VDD_XI10.XI24.MM17_s
+ N_VDD_XI10.XI24.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI10.XI27.MM17 N_XI10.XI27.NET31_XI10.XI27.MM17_d
+ N_XI10.XI27.NET27_XI10.XI27.MM17_g N_VDD_XI10.XI27.MM17_s
+ N_VDD_XI10.XI27.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI10.XI22.MM17 N_XI10.XI22.NET31_XI10.XI22.MM17_d
+ N_XI10.XI22.NET27_XI10.XI22.MM17_g N_VDD_XI10.XI22.MM17_s
+ N_VDD_XI10.XI22.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI10.XI21.MM17 N_XI10.XI21.NET31_XI10.XI21.MM17_d
+ N_XI10.XI21.NET27_XI10.XI21.MM17_g N_VDD_XI10.XI21.MM17_s
+ N_VDD_XI10.XI21.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI10.XI23.MM17 N_XI10.XI23.NET31_XI10.XI23.MM17_d
+ N_XI10.XI23.NET27_XI10.XI23.MM17_g N_VDD_XI10.XI23.MM17_s
+ N_VDD_XI10.XI23.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI10.XI19.MM17 N_XI10.XI19.NET31_XI10.XI19.MM17_d
+ N_XI10.XI19.NET27_XI10.XI19.MM17_g N_VDD_XI10.XI19.MM17_s
+ N_VDD_XI10.XI19.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI10.XI20.MM17 N_XI10.XI20.NET31_XI10.XI20.MM17_d
+ N_XI10.XI20.NET27_XI10.XI20.MM17_g N_VDD_XI10.XI20.MM17_s
+ N_VDD_XI10.XI20.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI10.XI18.MM17 N_XI10.XI18.NET31_XI10.XI18.MM17_d
+ N_XI10.XI18.NET27_XI10.XI18.MM17_g N_VDD_XI10.XI18.MM17_s
+ N_VDD_XI10.XI18.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI10.XI17.MM17 N_XI10.XI17.NET31_XI10.XI17.MM17_d
+ N_XI10.XI17.NET27_XI10.XI17.MM17_g N_VDD_XI10.XI17.MM17_s
+ N_VDD_XI10.XI17.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI10.XI0.MM37 N_XI10.XI0.NET15_XI10.XI0.MM37_d N_XI10.XI0.CLKB_XI10.XI0.MM37_g
+ N_XI10.XI0.NET14_XI10.XI0.MM37_s N_VDD_XI10.XI0.XI0.MM1_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.125e-12 AS=9.375e-13 PD=3e-06 PS=2.75e-06
mXI10.XI30.MM27 N_XI10.XI30.NET31_XI10.XI30.MM27_d
+ N_XI10.XI30.NET35_XI10.XI30.MM27_g N_XI10.XI30.NET58_XI10.XI30.MM27_s
+ N_VDD_XI10.XI30.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=1.125e-12 AS=9.375e-13
+ PD=3e-06 PS=2.75e-06
mXI10.XI29.MM27 N_XI10.XI29.NET31_XI10.XI29.MM27_d
+ N_XI10.XI29.NET35_XI10.XI29.MM27_g N_XI10.XI29.NET58_XI10.XI29.MM27_s
+ N_VDD_XI10.XI29.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=1.125e-12 AS=9.375e-13
+ PD=3e-06 PS=2.75e-06
mXI10.XI31.MM27 N_XI10.XI31.NET31_XI10.XI31.MM27_d
+ N_XI10.XI31.NET35_XI10.XI31.MM27_g N_XI10.XI31.NET58_XI10.XI31.MM27_s
+ N_VDD_XI10.XI31.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=1.125e-12 AS=9.375e-13
+ PD=3e-06 PS=2.75e-06
mXI10.XI28.MM27 N_XI10.XI28.NET31_XI10.XI28.MM27_d
+ N_XI10.XI28.NET35_XI10.XI28.MM27_g N_XI10.XI28.NET58_XI10.XI28.MM27_s
+ N_VDD_XI10.XI28.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=1.125e-12 AS=9.375e-13
+ PD=3e-06 PS=2.75e-06
mXI10.XI25.MM27 N_XI10.XI25.NET31_XI10.XI25.MM27_d
+ N_XI10.XI25.NET35_XI10.XI25.MM27_g N_XI10.XI25.NET58_XI10.XI25.MM27_s
+ N_VDD_XI10.XI25.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=1.125e-12 AS=9.375e-13
+ PD=3e-06 PS=2.75e-06
mXI10.XI26.MM27 N_XI10.XI26.NET31_XI10.XI26.MM27_d
+ N_XI10.XI26.NET35_XI10.XI26.MM27_g N_XI10.XI26.NET58_XI10.XI26.MM27_s
+ N_VDD_XI10.XI26.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=1.125e-12 AS=9.375e-13
+ PD=3e-06 PS=2.75e-06
mXI10.XI24.MM27 N_XI10.XI24.NET31_XI10.XI24.MM27_d
+ N_XI10.XI24.NET35_XI10.XI24.MM27_g N_XI10.XI24.NET58_XI10.XI24.MM27_s
+ N_VDD_XI10.XI24.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=1.125e-12 AS=9.375e-13
+ PD=3e-06 PS=2.75e-06
mXI10.XI27.MM27 N_XI10.XI27.NET31_XI10.XI27.MM27_d
+ N_XI10.XI27.NET35_XI10.XI27.MM27_g N_XI10.XI27.NET58_XI10.XI27.MM27_s
+ N_VDD_XI10.XI27.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=1.125e-12 AS=9.375e-13
+ PD=3e-06 PS=2.75e-06
mXI10.XI22.MM27 N_XI10.XI22.NET31_XI10.XI22.MM27_d
+ N_XI10.XI22.NET35_XI10.XI22.MM27_g N_XI10.XI22.NET58_XI10.XI22.MM27_s
+ N_VDD_XI10.XI22.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=1.125e-12 AS=9.375e-13
+ PD=3e-06 PS=2.75e-06
mXI10.XI21.MM27 N_XI10.XI21.NET31_XI10.XI21.MM27_d
+ N_XI10.XI21.NET35_XI10.XI21.MM27_g N_XI10.XI21.NET58_XI10.XI21.MM27_s
+ N_VDD_XI10.XI21.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=1.125e-12 AS=9.375e-13
+ PD=3e-06 PS=2.75e-06
mXI10.XI23.MM27 N_XI10.XI23.NET31_XI10.XI23.MM27_d
+ N_XI10.XI23.NET35_XI10.XI23.MM27_g N_XI10.XI23.NET58_XI10.XI23.MM27_s
+ N_VDD_XI10.XI23.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=1.125e-12 AS=9.375e-13
+ PD=3e-06 PS=2.75e-06
mXI10.XI19.MM27 N_XI10.XI19.NET31_XI10.XI19.MM27_d
+ N_XI10.XI19.NET35_XI10.XI19.MM27_g N_XI10.XI19.NET58_XI10.XI19.MM27_s
+ N_VDD_XI10.XI19.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=1.125e-12 AS=9.375e-13
+ PD=3e-06 PS=2.75e-06
mXI10.XI20.MM27 N_XI10.XI20.NET31_XI10.XI20.MM27_d
+ N_XI10.XI20.NET35_XI10.XI20.MM27_g N_XI10.XI20.NET58_XI10.XI20.MM27_s
+ N_VDD_XI10.XI20.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=1.125e-12 AS=9.375e-13
+ PD=3e-06 PS=2.75e-06
mXI10.XI18.MM27 N_XI10.XI18.NET31_XI10.XI18.MM27_d
+ N_XI10.XI18.NET35_XI10.XI18.MM27_g N_XI10.XI18.NET58_XI10.XI18.MM27_s
+ N_VDD_XI10.XI18.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=1.125e-12 AS=9.375e-13
+ PD=3e-06 PS=2.75e-06
mXI10.XI17.MM27 N_XI10.XI17.NET31_XI10.XI17.MM27_d
+ N_XI10.XI17.NET35_XI10.XI17.MM27_g N_XI10.XI17.NET58_XI10.XI17.MM27_s
+ N_VDD_XI10.XI17.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=1.125e-12 AS=9.375e-13
+ PD=3e-06 PS=2.75e-06
mXI10.XI0.MM13 N_NET256_XI10.XI0.MM13_d N_XI10.XI0.NET14_XI10.XI0.MM13_g
+ N_VDD_XI10.XI0.MM13_s N_VDD_XI10.XI0.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI10.XI30.MM3 N_XI10.XI30.NET15_XI10.XI30.MM3_d
+ N_XI10.XI30.NET58_XI10.XI30.MM3_g N_VDD_XI10.XI30.MM3_s
+ N_VDD_XI10.XI30.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI10.XI29.MM3 N_XI10.XI29.NET15_XI10.XI29.MM3_d
+ N_XI10.XI29.NET58_XI10.XI29.MM3_g N_VDD_XI10.XI29.MM3_s
+ N_VDD_XI10.XI29.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI10.XI31.MM3 N_XI10.XI31.NET15_XI10.XI31.MM3_d
+ N_XI10.XI31.NET58_XI10.XI31.MM3_g N_VDD_XI10.XI31.MM3_s
+ N_VDD_XI10.XI31.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI10.XI28.MM3 N_XI10.XI28.NET15_XI10.XI28.MM3_d
+ N_XI10.XI28.NET58_XI10.XI28.MM3_g N_VDD_XI10.XI28.MM3_s
+ N_VDD_XI10.XI28.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI10.XI25.MM3 N_XI10.XI25.NET15_XI10.XI25.MM3_d
+ N_XI10.XI25.NET58_XI10.XI25.MM3_g N_VDD_XI10.XI25.MM3_s
+ N_VDD_XI10.XI25.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI10.XI26.MM3 N_XI10.XI26.NET15_XI10.XI26.MM3_d
+ N_XI10.XI26.NET58_XI10.XI26.MM3_g N_VDD_XI10.XI26.MM3_s
+ N_VDD_XI10.XI26.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI10.XI24.MM3 N_XI10.XI24.NET15_XI10.XI24.MM3_d
+ N_XI10.XI24.NET58_XI10.XI24.MM3_g N_VDD_XI10.XI24.MM3_s
+ N_VDD_XI10.XI24.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI10.XI27.MM3 N_XI10.XI27.NET15_XI10.XI27.MM3_d
+ N_XI10.XI27.NET58_XI10.XI27.MM3_g N_VDD_XI10.XI27.MM3_s
+ N_VDD_XI10.XI27.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI10.XI22.MM3 N_XI10.XI22.NET15_XI10.XI22.MM3_d
+ N_XI10.XI22.NET58_XI10.XI22.MM3_g N_VDD_XI10.XI22.MM3_s
+ N_VDD_XI10.XI22.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI10.XI21.MM3 N_XI10.XI21.NET15_XI10.XI21.MM3_d
+ N_XI10.XI21.NET58_XI10.XI21.MM3_g N_VDD_XI10.XI21.MM3_s
+ N_VDD_XI10.XI21.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI10.XI23.MM3 N_XI10.XI23.NET15_XI10.XI23.MM3_d
+ N_XI10.XI23.NET58_XI10.XI23.MM3_g N_VDD_XI10.XI23.MM3_s
+ N_VDD_XI10.XI23.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI10.XI19.MM3 N_XI10.XI19.NET15_XI10.XI19.MM3_d
+ N_XI10.XI19.NET58_XI10.XI19.MM3_g N_VDD_XI10.XI19.MM3_s
+ N_VDD_XI10.XI19.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI10.XI20.MM3 N_XI10.XI20.NET15_XI10.XI20.MM3_d
+ N_XI10.XI20.NET58_XI10.XI20.MM3_g N_VDD_XI10.XI20.MM3_s
+ N_VDD_XI10.XI20.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI10.XI18.MM3 N_XI10.XI18.NET15_XI10.XI18.MM3_d
+ N_XI10.XI18.NET58_XI10.XI18.MM3_g N_VDD_XI10.XI18.MM3_s
+ N_VDD_XI10.XI18.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI10.XI17.MM3 N_XI10.XI17.NET15_XI10.XI17.MM3_d
+ N_XI10.XI17.NET58_XI10.XI17.MM3_g N_VDD_XI10.XI17.MM3_s
+ N_VDD_XI10.XI17.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI10.XI0.MM14 N_XI10.BAR_Q1_XI10.XI0.MM14_d N_NET256_XI10.XI0.MM14_g
+ N_VDD_XI10.XI0.MM14_s N_VDD_XI10.XI0.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI10.XI30.MM1 N_XI10.XI30.NET54_XI10.XI30.MM1_d
+ N_XI10.XI30.NET15_XI10.XI30.MM1_g N_VDD_XI10.XI30.MM1_s
+ N_VDD_XI10.XI30.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI10.XI29.MM1 N_XI10.XI29.NET54_XI10.XI29.MM1_d
+ N_XI10.XI29.NET15_XI10.XI29.MM1_g N_VDD_XI10.XI29.MM1_s
+ N_VDD_XI10.XI29.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI10.XI31.MM1 N_XI10.XI31.NET54_XI10.XI31.MM1_d
+ N_XI10.XI31.NET15_XI10.XI31.MM1_g N_VDD_XI10.XI31.MM1_s
+ N_VDD_XI10.XI31.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI10.XI28.MM1 N_XI10.XI28.NET54_XI10.XI28.MM1_d
+ N_XI10.XI28.NET15_XI10.XI28.MM1_g N_VDD_XI10.XI28.MM1_s
+ N_VDD_XI10.XI28.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI10.XI25.MM1 N_XI10.XI25.NET54_XI10.XI25.MM1_d
+ N_XI10.XI25.NET15_XI10.XI25.MM1_g N_VDD_XI10.XI25.MM1_s
+ N_VDD_XI10.XI25.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI10.XI26.MM1 N_XI10.XI26.NET54_XI10.XI26.MM1_d
+ N_XI10.XI26.NET15_XI10.XI26.MM1_g N_VDD_XI10.XI26.MM1_s
+ N_VDD_XI10.XI26.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI10.XI24.MM1 N_XI10.XI24.NET54_XI10.XI24.MM1_d
+ N_XI10.XI24.NET15_XI10.XI24.MM1_g N_VDD_XI10.XI24.MM1_s
+ N_VDD_XI10.XI24.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI10.XI27.MM1 N_XI10.XI27.NET54_XI10.XI27.MM1_d
+ N_XI10.XI27.NET15_XI10.XI27.MM1_g N_VDD_XI10.XI27.MM1_s
+ N_VDD_XI10.XI27.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI10.XI22.MM1 N_XI10.XI22.NET54_XI10.XI22.MM1_d
+ N_XI10.XI22.NET15_XI10.XI22.MM1_g N_VDD_XI10.XI22.MM1_s
+ N_VDD_XI10.XI22.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI10.XI21.MM1 N_XI10.XI21.NET54_XI10.XI21.MM1_d
+ N_XI10.XI21.NET15_XI10.XI21.MM1_g N_VDD_XI10.XI21.MM1_s
+ N_VDD_XI10.XI21.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI10.XI23.MM1 N_XI10.XI23.NET54_XI10.XI23.MM1_d
+ N_XI10.XI23.NET15_XI10.XI23.MM1_g N_VDD_XI10.XI23.MM1_s
+ N_VDD_XI10.XI23.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI10.XI19.MM1 N_XI10.XI19.NET54_XI10.XI19.MM1_d
+ N_XI10.XI19.NET15_XI10.XI19.MM1_g N_VDD_XI10.XI19.MM1_s
+ N_VDD_XI10.XI19.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI10.XI20.MM1 N_XI10.XI20.NET54_XI10.XI20.MM1_d
+ N_XI10.XI20.NET15_XI10.XI20.MM1_g N_VDD_XI10.XI20.MM1_s
+ N_VDD_XI10.XI20.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI10.XI18.MM1 N_XI10.XI18.NET54_XI10.XI18.MM1_d
+ N_XI10.XI18.NET15_XI10.XI18.MM1_g N_VDD_XI10.XI18.MM1_s
+ N_VDD_XI10.XI18.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI10.XI17.MM1 N_XI10.XI17.NET54_XI10.XI17.MM1_d
+ N_XI10.XI17.NET15_XI10.XI17.MM1_g N_VDD_XI10.XI17.MM1_s
+ N_VDD_XI10.XI17.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI10.XI0.MM39 N_XI10.XI0.NET14_XI10.XI0.MM39_d N_XI10.XI0.NET35_XI10.XI0.MM39_g
+ N_XI10.BAR_Q1_XI10.XI0.MM39_s N_VDD_XI10.XI0.XI0.MM1_b P_18 L=1.8e-07
+ W=1.5e-06 AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI10.XI30.MM35 N_XI10.XI30.NET58_XI10.XI30.MM35_d
+ N_XI10.XI30.CLKB_XI10.XI30.MM35_g N_XI10.XI30.NET54_XI10.XI30.MM35_s
+ N_VDD_XI10.XI30.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI10.XI29.MM35 N_XI10.XI29.NET58_XI10.XI29.MM35_d
+ N_XI10.XI29.CLKB_XI10.XI29.MM35_g N_XI10.XI29.NET54_XI10.XI29.MM35_s
+ N_VDD_XI10.XI29.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI10.XI31.MM35 N_XI10.XI31.NET58_XI10.XI31.MM35_d
+ N_XI10.XI31.CLKB_XI10.XI31.MM35_g N_XI10.XI31.NET54_XI10.XI31.MM35_s
+ N_VDD_XI10.XI31.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI10.XI28.MM35 N_XI10.XI28.NET58_XI10.XI28.MM35_d
+ N_XI10.XI28.CLKB_XI10.XI28.MM35_g N_XI10.XI28.NET54_XI10.XI28.MM35_s
+ N_VDD_XI10.XI28.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI10.XI25.MM35 N_XI10.XI25.NET58_XI10.XI25.MM35_d
+ N_XI10.XI25.CLKB_XI10.XI25.MM35_g N_XI10.XI25.NET54_XI10.XI25.MM35_s
+ N_VDD_XI10.XI25.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI10.XI26.MM35 N_XI10.XI26.NET58_XI10.XI26.MM35_d
+ N_XI10.XI26.CLKB_XI10.XI26.MM35_g N_XI10.XI26.NET54_XI10.XI26.MM35_s
+ N_VDD_XI10.XI26.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI10.XI24.MM35 N_XI10.XI24.NET58_XI10.XI24.MM35_d
+ N_XI10.XI24.CLKB_XI10.XI24.MM35_g N_XI10.XI24.NET54_XI10.XI24.MM35_s
+ N_VDD_XI10.XI24.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI10.XI27.MM35 N_XI10.XI27.NET58_XI10.XI27.MM35_d
+ N_XI10.XI27.CLKB_XI10.XI27.MM35_g N_XI10.XI27.NET54_XI10.XI27.MM35_s
+ N_VDD_XI10.XI27.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI10.XI22.MM35 N_XI10.XI22.NET58_XI10.XI22.MM35_d
+ N_XI10.XI22.CLKB_XI10.XI22.MM35_g N_XI10.XI22.NET54_XI10.XI22.MM35_s
+ N_VDD_XI10.XI22.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI10.XI21.MM35 N_XI10.XI21.NET58_XI10.XI21.MM35_d
+ N_XI10.XI21.CLKB_XI10.XI21.MM35_g N_XI10.XI21.NET54_XI10.XI21.MM35_s
+ N_VDD_XI10.XI21.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI10.XI23.MM35 N_XI10.XI23.NET58_XI10.XI23.MM35_d
+ N_XI10.XI23.CLKB_XI10.XI23.MM35_g N_XI10.XI23.NET54_XI10.XI23.MM35_s
+ N_VDD_XI10.XI23.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI10.XI19.MM35 N_XI10.XI19.NET58_XI10.XI19.MM35_d
+ N_XI10.XI19.CLKB_XI10.XI19.MM35_g N_XI10.XI19.NET54_XI10.XI19.MM35_s
+ N_VDD_XI10.XI19.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI10.XI20.MM35 N_XI10.XI20.NET58_XI10.XI20.MM35_d
+ N_XI10.XI20.CLKB_XI10.XI20.MM35_g N_XI10.XI20.NET54_XI10.XI20.MM35_s
+ N_VDD_XI10.XI20.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI10.XI18.MM35 N_XI10.XI18.NET58_XI10.XI18.MM35_d
+ N_XI10.XI18.CLKB_XI10.XI18.MM35_g N_XI10.XI18.NET54_XI10.XI18.MM35_s
+ N_VDD_XI10.XI18.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI10.XI17.MM35 N_XI10.XI17.NET58_XI10.XI17.MM35_d
+ N_XI10.XI17.CLKB_XI10.XI17.MM35_g N_XI10.XI17.NET54_XI10.XI17.MM35_s
+ N_VDD_XI10.XI17.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI10.XI30.MM37 N_XI10.XI30.NET15_XI10.XI30.MM37_d
+ N_XI10.XI30.CLKB_XI10.XI30.MM37_g N_XI10.XI30.NET14_XI10.XI30.MM37_s
+ N_VDD_XI10.XI30.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=1.125e-12 AS=9.375e-13
+ PD=3e-06 PS=2.75e-06
mXI10.XI29.MM37 N_XI10.XI29.NET15_XI10.XI29.MM37_d
+ N_XI10.XI29.CLKB_XI10.XI29.MM37_g N_XI10.XI29.NET14_XI10.XI29.MM37_s
+ N_VDD_XI10.XI29.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=1.125e-12 AS=9.375e-13
+ PD=3e-06 PS=2.75e-06
mXI10.XI31.MM37 N_XI10.XI31.NET15_XI10.XI31.MM37_d
+ N_XI10.XI31.CLKB_XI10.XI31.MM37_g N_XI10.XI31.NET14_XI10.XI31.MM37_s
+ N_VDD_XI10.XI31.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=1.125e-12 AS=9.375e-13
+ PD=3e-06 PS=2.75e-06
mXI10.XI28.MM37 N_XI10.XI28.NET15_XI10.XI28.MM37_d
+ N_XI10.XI28.CLKB_XI10.XI28.MM37_g N_XI10.XI28.NET14_XI10.XI28.MM37_s
+ N_VDD_XI10.XI28.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=1.125e-12 AS=9.375e-13
+ PD=3e-06 PS=2.75e-06
mXI10.XI25.MM37 N_XI10.XI25.NET15_XI10.XI25.MM37_d
+ N_XI10.XI25.CLKB_XI10.XI25.MM37_g N_XI10.XI25.NET14_XI10.XI25.MM37_s
+ N_VDD_XI10.XI25.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=1.125e-12 AS=9.375e-13
+ PD=3e-06 PS=2.75e-06
mXI10.XI26.MM37 N_XI10.XI26.NET15_XI10.XI26.MM37_d
+ N_XI10.XI26.CLKB_XI10.XI26.MM37_g N_XI10.XI26.NET14_XI10.XI26.MM37_s
+ N_VDD_XI10.XI26.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=1.125e-12 AS=9.375e-13
+ PD=3e-06 PS=2.75e-06
mXI10.XI24.MM37 N_XI10.XI24.NET15_XI10.XI24.MM37_d
+ N_XI10.XI24.CLKB_XI10.XI24.MM37_g N_XI10.XI24.NET14_XI10.XI24.MM37_s
+ N_VDD_XI10.XI24.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=1.125e-12 AS=9.375e-13
+ PD=3e-06 PS=2.75e-06
mXI10.XI27.MM37 N_XI10.XI27.NET15_XI10.XI27.MM37_d
+ N_XI10.XI27.CLKB_XI10.XI27.MM37_g N_XI10.XI27.NET14_XI10.XI27.MM37_s
+ N_VDD_XI10.XI27.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=1.125e-12 AS=9.375e-13
+ PD=3e-06 PS=2.75e-06
mXI10.XI22.MM37 N_XI10.XI22.NET15_XI10.XI22.MM37_d
+ N_XI10.XI22.CLKB_XI10.XI22.MM37_g N_XI10.XI22.NET14_XI10.XI22.MM37_s
+ N_VDD_XI10.XI22.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=1.125e-12 AS=9.375e-13
+ PD=3e-06 PS=2.75e-06
mXI10.XI21.MM37 N_XI10.XI21.NET15_XI10.XI21.MM37_d
+ N_XI10.XI21.CLKB_XI10.XI21.MM37_g N_XI10.XI21.NET14_XI10.XI21.MM37_s
+ N_VDD_XI10.XI21.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=1.125e-12 AS=9.375e-13
+ PD=3e-06 PS=2.75e-06
mXI10.XI23.MM37 N_XI10.XI23.NET15_XI10.XI23.MM37_d
+ N_XI10.XI23.CLKB_XI10.XI23.MM37_g N_XI10.XI23.NET14_XI10.XI23.MM37_s
+ N_VDD_XI10.XI23.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=1.125e-12 AS=9.375e-13
+ PD=3e-06 PS=2.75e-06
mXI10.XI19.MM37 N_XI10.XI19.NET15_XI10.XI19.MM37_d
+ N_XI10.XI19.CLKB_XI10.XI19.MM37_g N_XI10.XI19.NET14_XI10.XI19.MM37_s
+ N_VDD_XI10.XI19.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=1.125e-12 AS=9.375e-13
+ PD=3e-06 PS=2.75e-06
mXI10.XI20.MM37 N_XI10.XI20.NET15_XI10.XI20.MM37_d
+ N_XI10.XI20.CLKB_XI10.XI20.MM37_g N_XI10.XI20.NET14_XI10.XI20.MM37_s
+ N_VDD_XI10.XI20.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=1.125e-12 AS=9.375e-13
+ PD=3e-06 PS=2.75e-06
mXI10.XI18.MM37 N_XI10.XI18.NET15_XI10.XI18.MM37_d
+ N_XI10.XI18.CLKB_XI10.XI18.MM37_g N_XI10.XI18.NET14_XI10.XI18.MM37_s
+ N_VDD_XI10.XI18.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=1.125e-12 AS=9.375e-13
+ PD=3e-06 PS=2.75e-06
mXI10.XI17.MM37 N_XI10.XI17.NET15_XI10.XI17.MM37_d
+ N_XI10.XI17.CLKB_XI10.XI17.MM37_g N_XI10.XI17.NET14_XI10.XI17.MM37_s
+ N_VDD_XI10.XI17.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=1.125e-12 AS=9.375e-13
+ PD=3e-06 PS=2.75e-06
mXI9.XI97.XI4.MM1 N_XI9.XI97.NET39_XI9.XI97.XI4.MM1_d N_CIN1_XI9.XI97.XI4.MM1_g
+ N_VDD_XI9.XI97.XI4.MM1_s N_VDD_XI9.XI97.XI4.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI10.XI30.MM13 N_NET241_XI10.XI30.MM13_d N_XI10.XI30.NET14_XI10.XI30.MM13_g
+ N_VDD_XI10.XI30.MM13_s N_VDD_XI10.XI30.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI10.XI29.MM13 N_NET242_XI10.XI29.MM13_d N_XI10.XI29.NET14_XI10.XI29.MM13_g
+ N_VDD_XI10.XI29.MM13_s N_VDD_XI10.XI29.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI10.XI31.MM13 N_NET243_XI10.XI31.MM13_d N_XI10.XI31.NET14_XI10.XI31.MM13_g
+ N_VDD_XI10.XI31.MM13_s N_VDD_XI10.XI31.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI10.XI28.MM13 N_NET244_XI10.XI28.MM13_d N_XI10.XI28.NET14_XI10.XI28.MM13_g
+ N_VDD_XI10.XI28.MM13_s N_VDD_XI10.XI28.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI10.XI25.MM13 N_NET245_XI10.XI25.MM13_d N_XI10.XI25.NET14_XI10.XI25.MM13_g
+ N_VDD_XI10.XI25.MM13_s N_VDD_XI10.XI25.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI10.XI26.MM13 N_NET246_XI10.XI26.MM13_d N_XI10.XI26.NET14_XI10.XI26.MM13_g
+ N_VDD_XI10.XI26.MM13_s N_VDD_XI10.XI26.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI10.XI24.MM13 N_NET247_XI10.XI24.MM13_d N_XI10.XI24.NET14_XI10.XI24.MM13_g
+ N_VDD_XI10.XI24.MM13_s N_VDD_XI10.XI24.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI10.XI27.MM13 N_NET248_XI10.XI27.MM13_d N_XI10.XI27.NET14_XI10.XI27.MM13_g
+ N_VDD_XI10.XI27.MM13_s N_VDD_XI10.XI27.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI10.XI22.MM13 N_NET249_XI10.XI22.MM13_d N_XI10.XI22.NET14_XI10.XI22.MM13_g
+ N_VDD_XI10.XI22.MM13_s N_VDD_XI10.XI22.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI10.XI21.MM13 N_NET250_XI10.XI21.MM13_d N_XI10.XI21.NET14_XI10.XI21.MM13_g
+ N_VDD_XI10.XI21.MM13_s N_VDD_XI10.XI21.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI10.XI23.MM13 N_NET251_XI10.XI23.MM13_d N_XI10.XI23.NET14_XI10.XI23.MM13_g
+ N_VDD_XI10.XI23.MM13_s N_VDD_XI10.XI23.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI10.XI19.MM13 N_NET252_XI10.XI19.MM13_d N_XI10.XI19.NET14_XI10.XI19.MM13_g
+ N_VDD_XI10.XI19.MM13_s N_VDD_XI10.XI19.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI10.XI20.MM13 N_NET253_XI10.XI20.MM13_d N_XI10.XI20.NET14_XI10.XI20.MM13_g
+ N_VDD_XI10.XI20.MM13_s N_VDD_XI10.XI20.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI10.XI18.MM13 N_NET254_XI10.XI18.MM13_d N_XI10.XI18.NET14_XI10.XI18.MM13_g
+ N_VDD_XI10.XI18.MM13_s N_VDD_XI10.XI18.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI10.XI17.MM13 N_NET255_XI10.XI17.MM13_d N_XI10.XI17.NET14_XI10.XI17.MM13_g
+ N_VDD_XI10.XI17.MM13_s N_VDD_XI10.XI17.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI9.XI97.MM3 N_XI9.XI97.NET37_XI9.XI97.MM3_d N_XI9.XI97.NET39_XI9.XI97.MM3_g
+ N_VDD_XI9.XI97.MM3_s N_VDD_XI9.XI97.XI4.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=6.7125e-13 AS=9.675e-13 PD=8.95e-07 PS=2.79e-06
mXI9.XI97.MM1 N_NET192_XI9.XI97.MM1_d N_XI9.P1_XI9.XI97.MM1_g
+ N_XI9.XI97.NET37_XI9.XI97.MM1_s N_VDD_XI9.XI97.XI4.MM1_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.425e-12 AS=6.7125e-13 PD=1.9e-06 PS=8.95e-07
mXI10.XI30.MM14 N_XI10.BAR_Q16_XI10.XI30.MM14_d N_NET241_XI10.XI30.MM14_g
+ N_VDD_XI10.XI30.MM14_s N_VDD_XI10.XI30.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI10.XI29.MM14 N_XI10.BAR_Q15_XI10.XI29.MM14_d N_NET242_XI10.XI29.MM14_g
+ N_VDD_XI10.XI29.MM14_s N_VDD_XI10.XI29.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI10.XI31.MM14 N_XI10.BAR_Q14_XI10.XI31.MM14_d N_NET243_XI10.XI31.MM14_g
+ N_VDD_XI10.XI31.MM14_s N_VDD_XI10.XI31.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI10.XI28.MM14 N_XI10.BAR_Q13_XI10.XI28.MM14_d N_NET244_XI10.XI28.MM14_g
+ N_VDD_XI10.XI28.MM14_s N_VDD_XI10.XI28.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI10.XI25.MM14 N_XI10.BAR_Q12_XI10.XI25.MM14_d N_NET245_XI10.XI25.MM14_g
+ N_VDD_XI10.XI25.MM14_s N_VDD_XI10.XI25.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI10.XI26.MM14 N_XI10.BAR_Q11_XI10.XI26.MM14_d N_NET246_XI10.XI26.MM14_g
+ N_VDD_XI10.XI26.MM14_s N_VDD_XI10.XI26.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI10.XI24.MM14 N_XI10.BAR_Q10_XI10.XI24.MM14_d N_NET247_XI10.XI24.MM14_g
+ N_VDD_XI10.XI24.MM14_s N_VDD_XI10.XI24.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI10.XI27.MM14 N_XI10.BAR_Q9_XI10.XI27.MM14_d N_NET248_XI10.XI27.MM14_g
+ N_VDD_XI10.XI27.MM14_s N_VDD_XI10.XI27.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI10.XI22.MM14 N_XI10.BAR_Q8_XI10.XI22.MM14_d N_NET249_XI10.XI22.MM14_g
+ N_VDD_XI10.XI22.MM14_s N_VDD_XI10.XI22.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI10.XI21.MM14 N_XI10.BAR_Q7_XI10.XI21.MM14_d N_NET250_XI10.XI21.MM14_g
+ N_VDD_XI10.XI21.MM14_s N_VDD_XI10.XI21.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI10.XI23.MM14 N_XI10.BAR_Q6_XI10.XI23.MM14_d N_NET251_XI10.XI23.MM14_g
+ N_VDD_XI10.XI23.MM14_s N_VDD_XI10.XI23.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI10.XI19.MM14 N_XI10.BAR_Q5_XI10.XI19.MM14_d N_NET252_XI10.XI19.MM14_g
+ N_VDD_XI10.XI19.MM14_s N_VDD_XI10.XI19.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI10.XI20.MM14 N_XI10.BAR_Q4_XI10.XI20.MM14_d N_NET253_XI10.XI20.MM14_g
+ N_VDD_XI10.XI20.MM14_s N_VDD_XI10.XI20.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI10.XI18.MM14 N_XI10.BAR_Q3_XI10.XI18.MM14_d N_NET254_XI10.XI18.MM14_g
+ N_VDD_XI10.XI18.MM14_s N_VDD_XI10.XI18.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI10.XI17.MM14 N_XI10.BAR_Q2_XI10.XI17.MM14_d N_NET255_XI10.XI17.MM14_g
+ N_VDD_XI10.XI17.MM14_s N_VDD_XI10.XI17.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI9.XI97.MM5 N_NET192_XI9.XI97.MM5_d N_XI9.XI97.NET43_XI9.XI97.MM5_g
+ N_XI9.XI97.NET25_XI9.XI97.MM5_s N_VDD_XI9.XI97.XI4.MM1_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.425e-12 AS=5.4375e-13 PD=1.9e-06 PS=7.25e-07
mXI10.XI30.MM39 N_XI10.XI30.NET14_XI10.XI30.MM39_d
+ N_XI10.XI30.NET35_XI10.XI30.MM39_g N_XI10.BAR_Q16_XI10.XI30.MM39_s
+ N_VDD_XI10.XI30.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI10.XI29.MM39 N_XI10.XI29.NET14_XI10.XI29.MM39_d
+ N_XI10.XI29.NET35_XI10.XI29.MM39_g N_XI10.BAR_Q15_XI10.XI29.MM39_s
+ N_VDD_XI10.XI29.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI10.XI31.MM39 N_XI10.XI31.NET14_XI10.XI31.MM39_d
+ N_XI10.XI31.NET35_XI10.XI31.MM39_g N_XI10.BAR_Q14_XI10.XI31.MM39_s
+ N_VDD_XI10.XI31.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI10.XI28.MM39 N_XI10.XI28.NET14_XI10.XI28.MM39_d
+ N_XI10.XI28.NET35_XI10.XI28.MM39_g N_XI10.BAR_Q13_XI10.XI28.MM39_s
+ N_VDD_XI10.XI28.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI10.XI25.MM39 N_XI10.XI25.NET14_XI10.XI25.MM39_d
+ N_XI10.XI25.NET35_XI10.XI25.MM39_g N_XI10.BAR_Q12_XI10.XI25.MM39_s
+ N_VDD_XI10.XI25.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI10.XI26.MM39 N_XI10.XI26.NET14_XI10.XI26.MM39_d
+ N_XI10.XI26.NET35_XI10.XI26.MM39_g N_XI10.BAR_Q11_XI10.XI26.MM39_s
+ N_VDD_XI10.XI26.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI10.XI24.MM39 N_XI10.XI24.NET14_XI10.XI24.MM39_d
+ N_XI10.XI24.NET35_XI10.XI24.MM39_g N_XI10.BAR_Q10_XI10.XI24.MM39_s
+ N_VDD_XI10.XI24.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI10.XI27.MM39 N_XI10.XI27.NET14_XI10.XI27.MM39_d
+ N_XI10.XI27.NET35_XI10.XI27.MM39_g N_XI10.BAR_Q9_XI10.XI27.MM39_s
+ N_VDD_XI10.XI27.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI10.XI22.MM39 N_XI10.XI22.NET14_XI10.XI22.MM39_d
+ N_XI10.XI22.NET35_XI10.XI22.MM39_g N_XI10.BAR_Q8_XI10.XI22.MM39_s
+ N_VDD_XI10.XI22.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI10.XI21.MM39 N_XI10.XI21.NET14_XI10.XI21.MM39_d
+ N_XI10.XI21.NET35_XI10.XI21.MM39_g N_XI10.BAR_Q7_XI10.XI21.MM39_s
+ N_VDD_XI10.XI21.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI10.XI23.MM39 N_XI10.XI23.NET14_XI10.XI23.MM39_d
+ N_XI10.XI23.NET35_XI10.XI23.MM39_g N_XI10.BAR_Q6_XI10.XI23.MM39_s
+ N_VDD_XI10.XI23.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI10.XI19.MM39 N_XI10.XI19.NET14_XI10.XI19.MM39_d
+ N_XI10.XI19.NET35_XI10.XI19.MM39_g N_XI10.BAR_Q5_XI10.XI19.MM39_s
+ N_VDD_XI10.XI19.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI10.XI20.MM39 N_XI10.XI20.NET14_XI10.XI20.MM39_d
+ N_XI10.XI20.NET35_XI10.XI20.MM39_g N_XI10.BAR_Q4_XI10.XI20.MM39_s
+ N_VDD_XI10.XI20.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI10.XI18.MM39 N_XI10.XI18.NET14_XI10.XI18.MM39_d
+ N_XI10.XI18.NET35_XI10.XI18.MM39_g N_XI10.BAR_Q3_XI10.XI18.MM39_s
+ N_VDD_XI10.XI18.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI10.XI17.MM39 N_XI10.XI17.NET14_XI10.XI17.MM39_d
+ N_XI10.XI17.NET35_XI10.XI17.MM39_g N_XI10.BAR_Q2_XI10.XI17.MM39_s
+ N_VDD_XI10.XI17.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI9.XI97.MM4 N_XI9.XI97.NET25_XI9.XI97.MM4_d N_CIN1_XI9.XI97.MM4_g
+ N_VDD_XI9.XI97.MM4_s N_VDD_XI9.XI97.XI4.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=5.4375e-13 AS=7.65e-13 PD=7.25e-07 PS=2.52e-06
mXI9.XI97.XI9.MM1 N_XI9.XI97.NET43_XI9.XI97.XI9.MM1_d
+ N_XI9.P1_XI9.XI97.XI9.MM1_g N_VDD_XI9.XI97.XI9.MM1_s N_VDD_XI9.XI97.XI4.MM1_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9.XI153.XI1.MM1 N_XI9.XI153.NET6_XI9.XI153.XI1.MM1_d
+ N_NET242_XI9.XI153.XI1.MM1_g N_VDD_XI9.XI153.XI1.MM1_s
+ N_VDD_XI9.XI153.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.35e-13
+ PD=7.4e-07 PS=2.48e-06
mXI9.XI154.XI1.MM1 N_XI9.XI154.NET6_XI9.XI154.XI1.MM1_d
+ N_NET243_XI9.XI154.XI1.MM1_g N_VDD_XI9.XI154.XI1.MM1_s
+ N_VDD_XI9.XI154.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.35e-13
+ PD=7.4e-07 PS=2.48e-06
mXI9.XI157.XI1.MM1 N_XI9.XI157.NET6_XI9.XI157.XI1.MM1_d
+ N_NET244_XI9.XI157.XI1.MM1_g N_VDD_XI9.XI157.XI1.MM1_s
+ N_VDD_XI9.XI157.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.35e-13
+ PD=7.4e-07 PS=2.48e-06
mXI9.XI156.XI1.MM1 N_XI9.XI156.NET6_XI9.XI156.XI1.MM1_d
+ N_NET245_XI9.XI156.XI1.MM1_g N_VDD_XI9.XI156.XI1.MM1_s
+ N_VDD_XI9.XI156.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.35e-13
+ PD=7.4e-07 PS=2.48e-06
mXI9.XI155.XI1.MM1 N_XI9.XI155.NET6_XI9.XI155.XI1.MM1_d
+ N_NET246_XI9.XI155.XI1.MM1_g N_VDD_XI9.XI155.XI1.MM1_s
+ N_VDD_XI9.XI155.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.35e-13
+ PD=7.4e-07 PS=2.48e-06
mXI9.XI133.XI1.MM1 N_XI9.XI133.NET6_XI9.XI133.XI1.MM1_d
+ N_NET247_XI9.XI133.XI1.MM1_g N_VDD_XI9.XI133.XI1.MM1_s
+ N_VDD_XI9.XI133.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.35e-13
+ PD=7.4e-07 PS=2.48e-06
mXI9.XI132.XI1.MM1 N_XI9.XI132.NET6_XI9.XI132.XI1.MM1_d
+ N_NET248_XI9.XI132.XI1.MM1_g N_VDD_XI9.XI132.XI1.MM1_s
+ N_VDD_XI9.XI132.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.35e-13
+ PD=7.4e-07 PS=2.48e-06
mXI9.XI131.XI1.MM1 N_XI9.XI131.NET6_XI9.XI131.XI1.MM1_d
+ N_NET249_XI9.XI131.XI1.MM1_g N_VDD_XI9.XI131.XI1.MM1_s
+ N_VDD_XI9.XI131.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.35e-13
+ PD=7.4e-07 PS=2.48e-06
mXI9.XI111.XI1.MM1 N_XI9.XI111.NET6_XI9.XI111.XI1.MM1_d
+ N_NET250_XI9.XI111.XI1.MM1_g N_VDD_XI9.XI111.XI1.MM1_s
+ N_VDD_XI9.XI111.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.35e-13
+ PD=7.4e-07 PS=2.48e-06
mXI9.XI110.XI1.MM1 N_XI9.XI110.NET6_XI9.XI110.XI1.MM1_d
+ N_NET251_XI9.XI110.XI1.MM1_g N_VDD_XI9.XI110.XI1.MM1_s
+ N_VDD_XI9.XI110.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.35e-13
+ PD=7.4e-07 PS=2.48e-06
mXI9.XI103.XI1.MM1 N_XI9.XI103.NET6_XI9.XI103.XI1.MM1_d
+ N_NET252_XI9.XI103.XI1.MM1_g N_VDD_XI9.XI103.XI1.MM1_s
+ N_VDD_XI9.XI103.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.35e-13
+ PD=7.4e-07 PS=2.48e-06
mXI9.XI102.XI1.MM1 N_XI9.XI102.NET6_XI9.XI102.XI1.MM1_d
+ N_NET253_XI9.XI102.XI1.MM1_g N_VDD_XI9.XI102.XI1.MM1_s
+ N_VDD_XI9.XI102.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.35e-13
+ PD=7.4e-07 PS=2.48e-06
mXI9.XI88.XI1.MM1 N_XI9.XI88.NET6_XI9.XI88.XI1.MM1_d N_NET254_XI9.XI88.XI1.MM1_g
+ N_VDD_XI9.XI88.XI1.MM1_s N_VDD_XI9.XI88.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=5.55e-13 AS=7.35e-13 PD=7.4e-07 PS=2.48e-06
mXI9.XI82.XI1.MM1 N_XI9.XI82.NET6_XI9.XI82.XI1.MM1_d N_NET255_XI9.XI82.XI1.MM1_g
+ N_VDD_XI9.XI82.XI1.MM1_s N_VDD_XI9.XI82.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=5.55e-13 AS=7.35e-13 PD=7.4e-07 PS=2.48e-06
mXI9.XI10.XI1.MM1 N_XI9.XI10.NET6_XI9.XI10.XI1.MM1_d N_NET256_XI9.XI10.XI1.MM1_g
+ N_VDD_XI9.XI10.XI1.MM1_s N_VDD_XI9.XI97.XI4.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=5.55e-13 AS=7.35e-13 PD=7.4e-07 PS=2.48e-06
mXI9.XI153.XI1.MM3 N_XI9.XI153.NET6_XI9.XI153.XI1.MM3_d
+ N_ACC14_XI9.XI153.XI1.MM3_g N_VDD_XI9.XI153.XI1.MM3_s
+ N_VDD_XI9.XI153.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.65e-13
+ PD=7.4e-07 PS=2.52e-06
mXI9.XI154.XI1.MM3 N_XI9.XI154.NET6_XI9.XI154.XI1.MM3_d
+ N_ACC13_XI9.XI154.XI1.MM3_g N_VDD_XI9.XI154.XI1.MM3_s
+ N_VDD_XI9.XI154.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.65e-13
+ PD=7.4e-07 PS=2.52e-06
mXI9.XI157.XI1.MM3 N_XI9.XI157.NET6_XI9.XI157.XI1.MM3_d
+ N_ACC12_XI9.XI157.XI1.MM3_g N_VDD_XI9.XI157.XI1.MM3_s
+ N_VDD_XI9.XI157.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.65e-13
+ PD=7.4e-07 PS=2.52e-06
mXI9.XI156.XI1.MM3 N_XI9.XI156.NET6_XI9.XI156.XI1.MM3_d
+ N_ACC11_XI9.XI156.XI1.MM3_g N_VDD_XI9.XI156.XI1.MM3_s
+ N_VDD_XI9.XI156.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.65e-13
+ PD=7.4e-07 PS=2.52e-06
mXI9.XI155.XI1.MM3 N_XI9.XI155.NET6_XI9.XI155.XI1.MM3_d
+ N_ACC10_XI9.XI155.XI1.MM3_g N_VDD_XI9.XI155.XI1.MM3_s
+ N_VDD_XI9.XI155.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.65e-13
+ PD=7.4e-07 PS=2.52e-06
mXI9.XI133.XI1.MM3 N_XI9.XI133.NET6_XI9.XI133.XI1.MM3_d
+ N_ACC9_XI9.XI133.XI1.MM3_g N_VDD_XI9.XI133.XI1.MM3_s N_VDD_XI9.XI133.XI1.MM1_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.65e-13 PD=7.4e-07 PS=2.52e-06
mXI9.XI132.XI1.MM3 N_XI9.XI132.NET6_XI9.XI132.XI1.MM3_d
+ N_ACC8_XI9.XI132.XI1.MM3_g N_VDD_XI9.XI132.XI1.MM3_s N_VDD_XI9.XI132.XI1.MM1_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.65e-13 PD=7.4e-07 PS=2.52e-06
mXI9.XI131.XI1.MM3 N_XI9.XI131.NET6_XI9.XI131.XI1.MM3_d
+ N_ACC7_XI9.XI131.XI1.MM3_g N_VDD_XI9.XI131.XI1.MM3_s N_VDD_XI9.XI131.XI1.MM1_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.65e-13 PD=7.4e-07 PS=2.52e-06
mXI9.XI111.XI1.MM3 N_XI9.XI111.NET6_XI9.XI111.XI1.MM3_d
+ N_ACC6_XI9.XI111.XI1.MM3_g N_VDD_XI9.XI111.XI1.MM3_s N_VDD_XI9.XI111.XI1.MM1_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.65e-13 PD=7.4e-07 PS=2.52e-06
mXI9.XI110.XI1.MM3 N_XI9.XI110.NET6_XI9.XI110.XI1.MM3_d
+ N_ACC5_XI9.XI110.XI1.MM3_g N_VDD_XI9.XI110.XI1.MM3_s N_VDD_XI9.XI110.XI1.MM1_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.65e-13 PD=7.4e-07 PS=2.52e-06
mXI9.XI103.XI1.MM3 N_XI9.XI103.NET6_XI9.XI103.XI1.MM3_d
+ N_ACC4_XI9.XI103.XI1.MM3_g N_VDD_XI9.XI103.XI1.MM3_s N_VDD_XI9.XI103.XI1.MM1_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.65e-13 PD=7.4e-07 PS=2.52e-06
mXI9.XI102.XI1.MM3 N_XI9.XI102.NET6_XI9.XI102.XI1.MM3_d
+ N_ACC3_XI9.XI102.XI1.MM3_g N_VDD_XI9.XI102.XI1.MM3_s N_VDD_XI9.XI102.XI1.MM1_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.65e-13 PD=7.4e-07 PS=2.52e-06
mXI9.XI88.XI1.MM3 N_XI9.XI88.NET6_XI9.XI88.XI1.MM3_d N_ACC2_XI9.XI88.XI1.MM3_g
+ N_VDD_XI9.XI88.XI1.MM3_s N_VDD_XI9.XI88.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=5.55e-13 AS=7.65e-13 PD=7.4e-07 PS=2.52e-06
mXI9.XI82.XI1.MM3 N_XI9.XI82.NET6_XI9.XI82.XI1.MM3_d N_ACC1_XI9.XI82.XI1.MM3_g
+ N_VDD_XI9.XI82.XI1.MM3_s N_VDD_XI9.XI82.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=5.55e-13 AS=7.65e-13 PD=7.4e-07 PS=2.52e-06
mXI9.XI10.XI1.MM3 N_XI9.XI10.NET6_XI9.XI10.XI1.MM3_d N_ACC0_XI9.XI10.XI1.MM3_g
+ N_VDD_XI9.XI10.XI1.MM3_s N_VDD_XI9.XI97.XI4.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=5.55e-13 AS=7.65e-13 PD=7.4e-07 PS=2.52e-06
mXI9.XI134.XI4.MM1 N_XI9.XI134.NET39_XI9.XI134.XI4.MM1_d
+ N_NET241_XI9.XI134.XI4.MM1_g N_VDD_XI9.XI134.XI4.MM1_s
+ N_VDD_XI9.XI134.XI4.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI9.XI153.XI0.MM1 N_XI9.G15_XI9.XI153.XI0.MM1_d
+ N_XI9.XI153.NET6_XI9.XI153.XI0.MM1_g N_VDD_XI9.XI153.XI0.MM1_s
+ N_VDD_XI9.XI153.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI9.XI154.XI0.MM1 N_XI9.G14_XI9.XI154.XI0.MM1_d
+ N_XI9.XI154.NET6_XI9.XI154.XI0.MM1_g N_VDD_XI9.XI154.XI0.MM1_s
+ N_VDD_XI9.XI154.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI9.XI157.XI0.MM1 N_XI9.G13_XI9.XI157.XI0.MM1_d
+ N_XI9.XI157.NET6_XI9.XI157.XI0.MM1_g N_VDD_XI9.XI157.XI0.MM1_s
+ N_VDD_XI9.XI157.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI9.XI156.XI0.MM1 N_XI9.G12_XI9.XI156.XI0.MM1_d
+ N_XI9.XI156.NET6_XI9.XI156.XI0.MM1_g N_VDD_XI9.XI156.XI0.MM1_s
+ N_VDD_XI9.XI156.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI9.XI155.XI0.MM1 N_XI9.G11_XI9.XI155.XI0.MM1_d
+ N_XI9.XI155.NET6_XI9.XI155.XI0.MM1_g N_VDD_XI9.XI155.XI0.MM1_s
+ N_VDD_XI9.XI155.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI9.XI133.XI0.MM1 N_XI9.G10_XI9.XI133.XI0.MM1_d
+ N_XI9.XI133.NET6_XI9.XI133.XI0.MM1_g N_VDD_XI9.XI133.XI0.MM1_s
+ N_VDD_XI9.XI133.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI9.XI132.XI0.MM1 N_XI9.G9_XI9.XI132.XI0.MM1_d
+ N_XI9.XI132.NET6_XI9.XI132.XI0.MM1_g N_VDD_XI9.XI132.XI0.MM1_s
+ N_VDD_XI9.XI132.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI9.XI131.XI0.MM1 N_XI9.G8_XI9.XI131.XI0.MM1_d
+ N_XI9.XI131.NET6_XI9.XI131.XI0.MM1_g N_VDD_XI9.XI131.XI0.MM1_s
+ N_VDD_XI9.XI131.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI9.XI111.XI0.MM1 N_XI9.G7_XI9.XI111.XI0.MM1_d
+ N_XI9.XI111.NET6_XI9.XI111.XI0.MM1_g N_VDD_XI9.XI111.XI0.MM1_s
+ N_VDD_XI9.XI111.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI9.XI110.XI0.MM1 N_XI9.G6_XI9.XI110.XI0.MM1_d
+ N_XI9.XI110.NET6_XI9.XI110.XI0.MM1_g N_VDD_XI9.XI110.XI0.MM1_s
+ N_VDD_XI9.XI110.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI9.XI103.XI0.MM1 N_XI9.G5_XI9.XI103.XI0.MM1_d
+ N_XI9.XI103.NET6_XI9.XI103.XI0.MM1_g N_VDD_XI9.XI103.XI0.MM1_s
+ N_VDD_XI9.XI103.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI9.XI102.XI0.MM1 N_XI9.G4_XI9.XI102.XI0.MM1_d
+ N_XI9.XI102.NET6_XI9.XI102.XI0.MM1_g N_VDD_XI9.XI102.XI0.MM1_s
+ N_VDD_XI9.XI102.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI9.XI88.XI0.MM1 N_XI9.G3_XI9.XI88.XI0.MM1_d N_XI9.XI88.NET6_XI9.XI88.XI0.MM1_g
+ N_VDD_XI9.XI88.XI0.MM1_s N_VDD_XI9.XI88.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9.XI82.XI0.MM1 N_XI9.G2_XI9.XI82.XI0.MM1_d N_XI9.XI82.NET6_XI9.XI82.XI0.MM1_g
+ N_VDD_XI9.XI82.XI0.MM1_s N_VDD_XI9.XI82.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9.XI10.XI0.MM1 N_XI9.G1_XI9.XI10.XI0.MM1_d N_XI9.XI10.NET6_XI9.XI10.XI0.MM1_g
+ N_VDD_XI9.XI10.XI0.MM1_s N_VDD_XI9.XI97.XI4.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9.XI134.MM3 N_XI9.XI134.NET37_XI9.XI134.MM3_d
+ N_XI9.XI134.NET39_XI9.XI134.MM3_g N_VDD_XI9.XI134.MM3_s
+ N_VDD_XI9.XI134.XI4.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=6.7125e-13 AS=9.675e-13
+ PD=8.95e-07 PS=2.79e-06
mXI9.XI134.MM1 N_XI9.P16_XI9.XI134.MM1_d N_ACC15_XI9.XI134.MM1_g
+ N_XI9.XI134.NET37_XI9.XI134.MM1_s N_VDD_XI9.XI134.XI4.MM1_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.425e-12 AS=6.7125e-13 PD=1.9e-06 PS=8.95e-07
mXI9.XI137.XI4.MM1 N_XI9.XI137.NET39_XI9.XI137.XI4.MM1_d
+ N_NET242_XI9.XI137.XI4.MM1_g N_VDD_XI9.XI137.XI4.MM1_s
+ N_VDD_XI9.XI153.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI9.XI140.XI4.MM1 N_XI9.XI140.NET39_XI9.XI140.XI4.MM1_d
+ N_NET243_XI9.XI140.XI4.MM1_g N_VDD_XI9.XI140.XI4.MM1_s
+ N_VDD_XI9.XI154.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI9.XI149.XI4.MM1 N_XI9.XI149.NET39_XI9.XI149.XI4.MM1_d
+ N_NET244_XI9.XI149.XI4.MM1_g N_VDD_XI9.XI149.XI4.MM1_s
+ N_VDD_XI9.XI157.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI9.XI146.XI4.MM1 N_XI9.XI146.NET39_XI9.XI146.XI4.MM1_d
+ N_NET245_XI9.XI146.XI4.MM1_g N_VDD_XI9.XI146.XI4.MM1_s
+ N_VDD_XI9.XI156.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI9.XI143.XI4.MM1 N_XI9.XI143.NET39_XI9.XI143.XI4.MM1_d
+ N_NET246_XI9.XI143.XI4.MM1_g N_VDD_XI9.XI143.XI4.MM1_s
+ N_VDD_XI9.XI155.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI9.XI128.XI4.MM1 N_XI9.XI128.NET39_XI9.XI128.XI4.MM1_d
+ N_NET247_XI9.XI128.XI4.MM1_g N_VDD_XI9.XI128.XI4.MM1_s
+ N_VDD_XI9.XI133.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI9.XI125.XI4.MM1 N_XI9.XI125.NET39_XI9.XI125.XI4.MM1_d
+ N_NET248_XI9.XI125.XI4.MM1_g N_VDD_XI9.XI125.XI4.MM1_s
+ N_VDD_XI9.XI132.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI9.XI122.XI4.MM1 N_XI9.XI122.NET39_XI9.XI122.XI4.MM1_d
+ N_NET249_XI9.XI122.XI4.MM1_g N_VDD_XI9.XI122.XI4.MM1_s
+ N_VDD_XI9.XI131.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI9.XI114.XI4.MM1 N_XI9.XI114.NET39_XI9.XI114.XI4.MM1_d
+ N_NET250_XI9.XI114.XI4.MM1_g N_VDD_XI9.XI114.XI4.MM1_s
+ N_VDD_XI9.XI111.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI9.XI109.XI4.MM1 N_XI9.XI109.NET39_XI9.XI109.XI4.MM1_d
+ N_NET251_XI9.XI109.XI4.MM1_g N_VDD_XI9.XI109.XI4.MM1_s
+ N_VDD_XI9.XI110.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI9.XI106.XI4.MM1 N_XI9.XI106.NET39_XI9.XI106.XI4.MM1_d
+ N_NET252_XI9.XI106.XI4.MM1_g N_VDD_XI9.XI106.XI4.MM1_s
+ N_VDD_XI9.XI103.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI9.XI101.XI4.MM1 N_XI9.XI101.NET39_XI9.XI101.XI4.MM1_d
+ N_NET253_XI9.XI101.XI4.MM1_g N_VDD_XI9.XI101.XI4.MM1_s
+ N_VDD_XI9.XI102.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI9.XI86.XI4.MM1 N_XI9.XI86.NET39_XI9.XI86.XI4.MM1_d
+ N_NET254_XI9.XI86.XI4.MM1_g N_VDD_XI9.XI86.XI4.MM1_s N_VDD_XI9.XI88.XI1.MM1_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9.XI80.XI4.MM1 N_XI9.XI80.NET39_XI9.XI80.XI4.MM1_d
+ N_NET255_XI9.XI80.XI4.MM1_g N_VDD_XI9.XI80.XI4.MM1_s N_VDD_XI9.XI82.XI1.MM1_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9.XI26.XI4.MM1 N_XI9.XI26.NET39_XI9.XI26.XI4.MM1_d
+ N_NET256_XI9.XI26.XI4.MM1_g N_VDD_XI9.XI26.XI4.MM1_s N_VDD_XI9.XI97.XI4.MM1_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9.XI134.MM5 N_XI9.P16_XI9.XI134.MM5_d N_XI9.XI134.NET43_XI9.XI134.MM5_g
+ N_XI9.XI134.NET25_XI9.XI134.MM5_s N_VDD_XI9.XI134.XI4.MM1_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.425e-12 AS=5.4375e-13 PD=1.9e-06 PS=7.25e-07
mXI9.XI137.MM3 N_XI9.XI137.NET37_XI9.XI137.MM3_d
+ N_XI9.XI137.NET39_XI9.XI137.MM3_g N_VDD_XI9.XI137.MM3_s
+ N_VDD_XI9.XI153.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=6.7125e-13 AS=9.675e-13
+ PD=8.95e-07 PS=2.79e-06
mXI9.XI140.MM3 N_XI9.XI140.NET37_XI9.XI140.MM3_d
+ N_XI9.XI140.NET39_XI9.XI140.MM3_g N_VDD_XI9.XI140.MM3_s
+ N_VDD_XI9.XI154.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=6.7125e-13 AS=9.675e-13
+ PD=8.95e-07 PS=2.79e-06
mXI9.XI149.MM3 N_XI9.XI149.NET37_XI9.XI149.MM3_d
+ N_XI9.XI149.NET39_XI9.XI149.MM3_g N_VDD_XI9.XI149.MM3_s
+ N_VDD_XI9.XI157.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=6.7125e-13 AS=9.675e-13
+ PD=8.95e-07 PS=2.79e-06
mXI9.XI146.MM3 N_XI9.XI146.NET37_XI9.XI146.MM3_d
+ N_XI9.XI146.NET39_XI9.XI146.MM3_g N_VDD_XI9.XI146.MM3_s
+ N_VDD_XI9.XI156.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=6.7125e-13 AS=9.675e-13
+ PD=8.95e-07 PS=2.79e-06
mXI9.XI143.MM3 N_XI9.XI143.NET37_XI9.XI143.MM3_d
+ N_XI9.XI143.NET39_XI9.XI143.MM3_g N_VDD_XI9.XI143.MM3_s
+ N_VDD_XI9.XI155.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=6.7125e-13 AS=9.675e-13
+ PD=8.95e-07 PS=2.79e-06
mXI9.XI128.MM3 N_XI9.XI128.NET37_XI9.XI128.MM3_d
+ N_XI9.XI128.NET39_XI9.XI128.MM3_g N_VDD_XI9.XI128.MM3_s
+ N_VDD_XI9.XI133.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=6.7125e-13 AS=9.675e-13
+ PD=8.95e-07 PS=2.79e-06
mXI9.XI125.MM3 N_XI9.XI125.NET37_XI9.XI125.MM3_d
+ N_XI9.XI125.NET39_XI9.XI125.MM3_g N_VDD_XI9.XI125.MM3_s
+ N_VDD_XI9.XI132.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=6.7125e-13 AS=9.675e-13
+ PD=8.95e-07 PS=2.79e-06
mXI9.XI122.MM3 N_XI9.XI122.NET37_XI9.XI122.MM3_d
+ N_XI9.XI122.NET39_XI9.XI122.MM3_g N_VDD_XI9.XI122.MM3_s
+ N_VDD_XI9.XI131.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=6.7125e-13 AS=9.675e-13
+ PD=8.95e-07 PS=2.79e-06
mXI9.XI114.MM3 N_XI9.XI114.NET37_XI9.XI114.MM3_d
+ N_XI9.XI114.NET39_XI9.XI114.MM3_g N_VDD_XI9.XI114.MM3_s
+ N_VDD_XI9.XI111.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=6.7125e-13 AS=9.675e-13
+ PD=8.95e-07 PS=2.79e-06
mXI9.XI109.MM3 N_XI9.XI109.NET37_XI9.XI109.MM3_d
+ N_XI9.XI109.NET39_XI9.XI109.MM3_g N_VDD_XI9.XI109.MM3_s
+ N_VDD_XI9.XI110.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=6.7125e-13 AS=9.675e-13
+ PD=8.95e-07 PS=2.79e-06
mXI9.XI106.MM3 N_XI9.XI106.NET37_XI9.XI106.MM3_d
+ N_XI9.XI106.NET39_XI9.XI106.MM3_g N_VDD_XI9.XI106.MM3_s
+ N_VDD_XI9.XI103.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=6.7125e-13 AS=9.675e-13
+ PD=8.95e-07 PS=2.79e-06
mXI9.XI101.MM3 N_XI9.XI101.NET37_XI9.XI101.MM3_d
+ N_XI9.XI101.NET39_XI9.XI101.MM3_g N_VDD_XI9.XI101.MM3_s
+ N_VDD_XI9.XI102.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=6.7125e-13 AS=9.675e-13
+ PD=8.95e-07 PS=2.79e-06
mXI9.XI86.MM3 N_XI9.XI86.NET37_XI9.XI86.MM3_d N_XI9.XI86.NET39_XI9.XI86.MM3_g
+ N_VDD_XI9.XI86.MM3_s N_VDD_XI9.XI88.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=6.7125e-13 AS=9.675e-13 PD=8.95e-07 PS=2.79e-06
mXI9.XI80.MM3 N_XI9.XI80.NET37_XI9.XI80.MM3_d N_XI9.XI80.NET39_XI9.XI80.MM3_g
+ N_VDD_XI9.XI80.MM3_s N_VDD_XI9.XI82.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=6.7125e-13 AS=9.675e-13 PD=8.95e-07 PS=2.79e-06
mXI9.XI26.MM3 N_XI9.XI26.NET37_XI9.XI26.MM3_d N_XI9.XI26.NET39_XI9.XI26.MM3_g
+ N_VDD_XI9.XI26.MM3_s N_VDD_XI9.XI97.XI4.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=6.7125e-13 AS=9.675e-13 PD=8.95e-07 PS=2.79e-06
mXI9.XI134.MM4 N_XI9.XI134.NET25_XI9.XI134.MM4_d N_NET241_XI9.XI134.MM4_g
+ N_VDD_XI9.XI134.MM4_s N_VDD_XI9.XI134.XI4.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=5.4375e-13 AS=7.65e-13 PD=7.25e-07 PS=2.52e-06
mXI9.XI137.MM1 N_XI9.P15_XI9.XI137.MM1_d N_ACC14_XI9.XI137.MM1_g
+ N_XI9.XI137.NET37_XI9.XI137.MM1_s N_VDD_XI9.XI153.XI1.MM1_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.425e-12 AS=6.7125e-13 PD=1.9e-06 PS=8.95e-07
mXI9.XI140.MM1 N_XI9.P14_XI9.XI140.MM1_d N_ACC13_XI9.XI140.MM1_g
+ N_XI9.XI140.NET37_XI9.XI140.MM1_s N_VDD_XI9.XI154.XI1.MM1_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.425e-12 AS=6.7125e-13 PD=1.9e-06 PS=8.95e-07
mXI9.XI149.MM1 N_XI9.P13_XI9.XI149.MM1_d N_ACC12_XI9.XI149.MM1_g
+ N_XI9.XI149.NET37_XI9.XI149.MM1_s N_VDD_XI9.XI157.XI1.MM1_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.425e-12 AS=6.7125e-13 PD=1.9e-06 PS=8.95e-07
mXI9.XI146.MM1 N_XI9.P12_XI9.XI146.MM1_d N_ACC11_XI9.XI146.MM1_g
+ N_XI9.XI146.NET37_XI9.XI146.MM1_s N_VDD_XI9.XI156.XI1.MM1_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.425e-12 AS=6.7125e-13 PD=1.9e-06 PS=8.95e-07
mXI9.XI143.MM1 N_XI9.P11_XI9.XI143.MM1_d N_ACC10_XI9.XI143.MM1_g
+ N_XI9.XI143.NET37_XI9.XI143.MM1_s N_VDD_XI9.XI155.XI1.MM1_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.425e-12 AS=6.7125e-13 PD=1.9e-06 PS=8.95e-07
mXI9.XI128.MM1 N_XI9.P10_XI9.XI128.MM1_d N_ACC9_XI9.XI128.MM1_g
+ N_XI9.XI128.NET37_XI9.XI128.MM1_s N_VDD_XI9.XI133.XI1.MM1_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.425e-12 AS=6.7125e-13 PD=1.9e-06 PS=8.95e-07
mXI9.XI125.MM1 N_XI9.P9_XI9.XI125.MM1_d N_ACC8_XI9.XI125.MM1_g
+ N_XI9.XI125.NET37_XI9.XI125.MM1_s N_VDD_XI9.XI132.XI1.MM1_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.425e-12 AS=6.7125e-13 PD=1.9e-06 PS=8.95e-07
mXI9.XI122.MM1 N_XI9.P8_XI9.XI122.MM1_d N_ACC7_XI9.XI122.MM1_g
+ N_XI9.XI122.NET37_XI9.XI122.MM1_s N_VDD_XI9.XI131.XI1.MM1_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.425e-12 AS=6.7125e-13 PD=1.9e-06 PS=8.95e-07
mXI9.XI114.MM1 N_XI9.P7_XI9.XI114.MM1_d N_ACC6_XI9.XI114.MM1_g
+ N_XI9.XI114.NET37_XI9.XI114.MM1_s N_VDD_XI9.XI111.XI1.MM1_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.425e-12 AS=6.7125e-13 PD=1.9e-06 PS=8.95e-07
mXI9.XI109.MM1 N_XI9.P6_XI9.XI109.MM1_d N_ACC5_XI9.XI109.MM1_g
+ N_XI9.XI109.NET37_XI9.XI109.MM1_s N_VDD_XI9.XI110.XI1.MM1_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.425e-12 AS=6.7125e-13 PD=1.9e-06 PS=8.95e-07
mXI9.XI106.MM1 N_XI9.P5_XI9.XI106.MM1_d N_ACC4_XI9.XI106.MM1_g
+ N_XI9.XI106.NET37_XI9.XI106.MM1_s N_VDD_XI9.XI103.XI1.MM1_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.425e-12 AS=6.7125e-13 PD=1.9e-06 PS=8.95e-07
mXI9.XI101.MM1 N_XI9.P4_XI9.XI101.MM1_d N_ACC3_XI9.XI101.MM1_g
+ N_XI9.XI101.NET37_XI9.XI101.MM1_s N_VDD_XI9.XI102.XI1.MM1_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.425e-12 AS=6.7125e-13 PD=1.9e-06 PS=8.95e-07
mXI9.XI86.MM1 N_XI9.P3_XI9.XI86.MM1_d N_ACC2_XI9.XI86.MM1_g
+ N_XI9.XI86.NET37_XI9.XI86.MM1_s N_VDD_XI9.XI88.XI1.MM1_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.425e-12 AS=6.7125e-13 PD=1.9e-06 PS=8.95e-07
mXI9.XI80.MM1 N_XI9.P2_XI9.XI80.MM1_d N_ACC1_XI9.XI80.MM1_g
+ N_XI9.XI80.NET37_XI9.XI80.MM1_s N_VDD_XI9.XI82.XI1.MM1_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.425e-12 AS=6.7125e-13 PD=1.9e-06 PS=8.95e-07
mXI9.XI26.MM1 N_XI9.P1_XI9.XI26.MM1_d N_ACC0_XI9.XI26.MM1_g
+ N_XI9.XI26.NET37_XI9.XI26.MM1_s N_VDD_XI9.XI97.XI4.MM1_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.425e-12 AS=6.7125e-13 PD=1.9e-06 PS=8.95e-07
mXI9.XI134.XI9.MM1 N_XI9.XI134.NET43_XI9.XI134.XI9.MM1_d
+ N_ACC15_XI9.XI134.XI9.MM1_g N_VDD_XI9.XI134.XI9.MM1_s
+ N_VDD_XI9.XI134.XI4.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI9.XI137.MM5 N_XI9.P15_XI9.XI137.MM5_d N_XI9.XI137.NET43_XI9.XI137.MM5_g
+ N_XI9.XI137.NET25_XI9.XI137.MM5_s N_VDD_XI9.XI153.XI1.MM1_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.425e-12 AS=5.4375e-13 PD=1.9e-06 PS=7.25e-07
mXI9.XI140.MM5 N_XI9.P14_XI9.XI140.MM5_d N_XI9.XI140.NET43_XI9.XI140.MM5_g
+ N_XI9.XI140.NET25_XI9.XI140.MM5_s N_VDD_XI9.XI154.XI1.MM1_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.425e-12 AS=5.4375e-13 PD=1.9e-06 PS=7.25e-07
mXI9.XI149.MM5 N_XI9.P13_XI9.XI149.MM5_d N_XI9.XI149.NET43_XI9.XI149.MM5_g
+ N_XI9.XI149.NET25_XI9.XI149.MM5_s N_VDD_XI9.XI157.XI1.MM1_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.425e-12 AS=5.4375e-13 PD=1.9e-06 PS=7.25e-07
mXI9.XI146.MM5 N_XI9.P12_XI9.XI146.MM5_d N_XI9.XI146.NET43_XI9.XI146.MM5_g
+ N_XI9.XI146.NET25_XI9.XI146.MM5_s N_VDD_XI9.XI156.XI1.MM1_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.425e-12 AS=5.4375e-13 PD=1.9e-06 PS=7.25e-07
mXI9.XI143.MM5 N_XI9.P11_XI9.XI143.MM5_d N_XI9.XI143.NET43_XI9.XI143.MM5_g
+ N_XI9.XI143.NET25_XI9.XI143.MM5_s N_VDD_XI9.XI155.XI1.MM1_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.425e-12 AS=5.4375e-13 PD=1.9e-06 PS=7.25e-07
mXI9.XI128.MM5 N_XI9.P10_XI9.XI128.MM5_d N_XI9.XI128.NET43_XI9.XI128.MM5_g
+ N_XI9.XI128.NET25_XI9.XI128.MM5_s N_VDD_XI9.XI133.XI1.MM1_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.425e-12 AS=5.4375e-13 PD=1.9e-06 PS=7.25e-07
mXI9.XI125.MM5 N_XI9.P9_XI9.XI125.MM5_d N_XI9.XI125.NET43_XI9.XI125.MM5_g
+ N_XI9.XI125.NET25_XI9.XI125.MM5_s N_VDD_XI9.XI132.XI1.MM1_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.425e-12 AS=5.4375e-13 PD=1.9e-06 PS=7.25e-07
mXI9.XI122.MM5 N_XI9.P8_XI9.XI122.MM5_d N_XI9.XI122.NET43_XI9.XI122.MM5_g
+ N_XI9.XI122.NET25_XI9.XI122.MM5_s N_VDD_XI9.XI131.XI1.MM1_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.425e-12 AS=5.4375e-13 PD=1.9e-06 PS=7.25e-07
mXI9.XI114.MM5 N_XI9.P7_XI9.XI114.MM5_d N_XI9.XI114.NET43_XI9.XI114.MM5_g
+ N_XI9.XI114.NET25_XI9.XI114.MM5_s N_VDD_XI9.XI111.XI1.MM1_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.425e-12 AS=5.4375e-13 PD=1.9e-06 PS=7.25e-07
mXI9.XI109.MM5 N_XI9.P6_XI9.XI109.MM5_d N_XI9.XI109.NET43_XI9.XI109.MM5_g
+ N_XI9.XI109.NET25_XI9.XI109.MM5_s N_VDD_XI9.XI110.XI1.MM1_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.425e-12 AS=5.4375e-13 PD=1.9e-06 PS=7.25e-07
mXI9.XI106.MM5 N_XI9.P5_XI9.XI106.MM5_d N_XI9.XI106.NET43_XI9.XI106.MM5_g
+ N_XI9.XI106.NET25_XI9.XI106.MM5_s N_VDD_XI9.XI103.XI1.MM1_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.425e-12 AS=5.4375e-13 PD=1.9e-06 PS=7.25e-07
mXI9.XI101.MM5 N_XI9.P4_XI9.XI101.MM5_d N_XI9.XI101.NET43_XI9.XI101.MM5_g
+ N_XI9.XI101.NET25_XI9.XI101.MM5_s N_VDD_XI9.XI102.XI1.MM1_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.425e-12 AS=5.4375e-13 PD=1.9e-06 PS=7.25e-07
mXI9.XI86.MM5 N_XI9.P3_XI9.XI86.MM5_d N_XI9.XI86.NET43_XI9.XI86.MM5_g
+ N_XI9.XI86.NET25_XI9.XI86.MM5_s N_VDD_XI9.XI88.XI1.MM1_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.425e-12 AS=5.4375e-13 PD=1.9e-06 PS=7.25e-07
mXI9.XI80.MM5 N_XI9.P2_XI9.XI80.MM5_d N_XI9.XI80.NET43_XI9.XI80.MM5_g
+ N_XI9.XI80.NET25_XI9.XI80.MM5_s N_VDD_XI9.XI82.XI1.MM1_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.425e-12 AS=5.4375e-13 PD=1.9e-06 PS=7.25e-07
mXI9.XI26.MM5 N_XI9.P1_XI9.XI26.MM5_d N_XI9.XI26.NET43_XI9.XI26.MM5_g
+ N_XI9.XI26.NET25_XI9.XI26.MM5_s N_VDD_XI9.XI97.XI4.MM1_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.425e-12 AS=5.4375e-13 PD=1.9e-06 PS=7.25e-07
mXI9.XI137.MM4 N_XI9.XI137.NET25_XI9.XI137.MM4_d N_NET242_XI9.XI137.MM4_g
+ N_VDD_XI9.XI137.MM4_s N_VDD_XI9.XI153.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=5.4375e-13 AS=7.65e-13 PD=7.25e-07 PS=2.52e-06
mXI9.XI140.MM4 N_XI9.XI140.NET25_XI9.XI140.MM4_d N_NET243_XI9.XI140.MM4_g
+ N_VDD_XI9.XI140.MM4_s N_VDD_XI9.XI154.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=5.4375e-13 AS=7.65e-13 PD=7.25e-07 PS=2.52e-06
mXI9.XI149.MM4 N_XI9.XI149.NET25_XI9.XI149.MM4_d N_NET244_XI9.XI149.MM4_g
+ N_VDD_XI9.XI149.MM4_s N_VDD_XI9.XI157.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=5.4375e-13 AS=7.65e-13 PD=7.25e-07 PS=2.52e-06
mXI9.XI146.MM4 N_XI9.XI146.NET25_XI9.XI146.MM4_d N_NET245_XI9.XI146.MM4_g
+ N_VDD_XI9.XI146.MM4_s N_VDD_XI9.XI156.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=5.4375e-13 AS=7.65e-13 PD=7.25e-07 PS=2.52e-06
mXI9.XI143.MM4 N_XI9.XI143.NET25_XI9.XI143.MM4_d N_NET246_XI9.XI143.MM4_g
+ N_VDD_XI9.XI143.MM4_s N_VDD_XI9.XI155.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=5.4375e-13 AS=7.65e-13 PD=7.25e-07 PS=2.52e-06
mXI9.XI128.MM4 N_XI9.XI128.NET25_XI9.XI128.MM4_d N_NET247_XI9.XI128.MM4_g
+ N_VDD_XI9.XI128.MM4_s N_VDD_XI9.XI133.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=5.4375e-13 AS=7.65e-13 PD=7.25e-07 PS=2.52e-06
mXI9.XI125.MM4 N_XI9.XI125.NET25_XI9.XI125.MM4_d N_NET248_XI9.XI125.MM4_g
+ N_VDD_XI9.XI125.MM4_s N_VDD_XI9.XI132.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=5.4375e-13 AS=7.65e-13 PD=7.25e-07 PS=2.52e-06
mXI9.XI122.MM4 N_XI9.XI122.NET25_XI9.XI122.MM4_d N_NET249_XI9.XI122.MM4_g
+ N_VDD_XI9.XI122.MM4_s N_VDD_XI9.XI131.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=5.4375e-13 AS=7.65e-13 PD=7.25e-07 PS=2.52e-06
mXI9.XI114.MM4 N_XI9.XI114.NET25_XI9.XI114.MM4_d N_NET250_XI9.XI114.MM4_g
+ N_VDD_XI9.XI114.MM4_s N_VDD_XI9.XI111.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=5.4375e-13 AS=7.65e-13 PD=7.25e-07 PS=2.52e-06
mXI9.XI109.MM4 N_XI9.XI109.NET25_XI9.XI109.MM4_d N_NET251_XI9.XI109.MM4_g
+ N_VDD_XI9.XI109.MM4_s N_VDD_XI9.XI110.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=5.4375e-13 AS=7.65e-13 PD=7.25e-07 PS=2.52e-06
mXI9.XI106.MM4 N_XI9.XI106.NET25_XI9.XI106.MM4_d N_NET252_XI9.XI106.MM4_g
+ N_VDD_XI9.XI106.MM4_s N_VDD_XI9.XI103.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=5.4375e-13 AS=7.65e-13 PD=7.25e-07 PS=2.52e-06
mXI9.XI101.MM4 N_XI9.XI101.NET25_XI9.XI101.MM4_d N_NET253_XI9.XI101.MM4_g
+ N_VDD_XI9.XI101.MM4_s N_VDD_XI9.XI102.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=5.4375e-13 AS=7.65e-13 PD=7.25e-07 PS=2.52e-06
mXI9.XI86.MM4 N_XI9.XI86.NET25_XI9.XI86.MM4_d N_NET254_XI9.XI86.MM4_g
+ N_VDD_XI9.XI86.MM4_s N_VDD_XI9.XI88.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=5.4375e-13 AS=7.65e-13 PD=7.25e-07 PS=2.52e-06
mXI9.XI80.MM4 N_XI9.XI80.NET25_XI9.XI80.MM4_d N_NET255_XI9.XI80.MM4_g
+ N_VDD_XI9.XI80.MM4_s N_VDD_XI9.XI82.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=5.4375e-13 AS=7.65e-13 PD=7.25e-07 PS=2.52e-06
mXI9.XI26.MM4 N_XI9.XI26.NET25_XI9.XI26.MM4_d N_NET256_XI9.XI26.MM4_g
+ N_VDD_XI9.XI26.MM4_s N_VDD_XI9.XI97.XI4.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=5.4375e-13 AS=7.65e-13 PD=7.25e-07 PS=2.52e-06
mXI9.XI137.XI9.MM1 N_XI9.XI137.NET43_XI9.XI137.XI9.MM1_d
+ N_ACC14_XI9.XI137.XI9.MM1_g N_VDD_XI9.XI137.XI9.MM1_s
+ N_VDD_XI9.XI153.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI9.XI140.XI9.MM1 N_XI9.XI140.NET43_XI9.XI140.XI9.MM1_d
+ N_ACC13_XI9.XI140.XI9.MM1_g N_VDD_XI9.XI140.XI9.MM1_s
+ N_VDD_XI9.XI154.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI9.XI149.XI9.MM1 N_XI9.XI149.NET43_XI9.XI149.XI9.MM1_d
+ N_ACC12_XI9.XI149.XI9.MM1_g N_VDD_XI9.XI149.XI9.MM1_s
+ N_VDD_XI9.XI157.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI9.XI146.XI9.MM1 N_XI9.XI146.NET43_XI9.XI146.XI9.MM1_d
+ N_ACC11_XI9.XI146.XI9.MM1_g N_VDD_XI9.XI146.XI9.MM1_s
+ N_VDD_XI9.XI156.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI9.XI143.XI9.MM1 N_XI9.XI143.NET43_XI9.XI143.XI9.MM1_d
+ N_ACC10_XI9.XI143.XI9.MM1_g N_VDD_XI9.XI143.XI9.MM1_s
+ N_VDD_XI9.XI155.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI9.XI128.XI9.MM1 N_XI9.XI128.NET43_XI9.XI128.XI9.MM1_d
+ N_ACC9_XI9.XI128.XI9.MM1_g N_VDD_XI9.XI128.XI9.MM1_s N_VDD_XI9.XI133.XI1.MM1_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9.XI125.XI9.MM1 N_XI9.XI125.NET43_XI9.XI125.XI9.MM1_d
+ N_ACC8_XI9.XI125.XI9.MM1_g N_VDD_XI9.XI125.XI9.MM1_s N_VDD_XI9.XI132.XI1.MM1_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9.XI122.XI9.MM1 N_XI9.XI122.NET43_XI9.XI122.XI9.MM1_d
+ N_ACC7_XI9.XI122.XI9.MM1_g N_VDD_XI9.XI122.XI9.MM1_s N_VDD_XI9.XI131.XI1.MM1_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9.XI114.XI9.MM1 N_XI9.XI114.NET43_XI9.XI114.XI9.MM1_d
+ N_ACC6_XI9.XI114.XI9.MM1_g N_VDD_XI9.XI114.XI9.MM1_s N_VDD_XI9.XI111.XI1.MM1_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9.XI109.XI9.MM1 N_XI9.XI109.NET43_XI9.XI109.XI9.MM1_d
+ N_ACC5_XI9.XI109.XI9.MM1_g N_VDD_XI9.XI109.XI9.MM1_s N_VDD_XI9.XI110.XI1.MM1_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9.XI106.XI9.MM1 N_XI9.XI106.NET43_XI9.XI106.XI9.MM1_d
+ N_ACC4_XI9.XI106.XI9.MM1_g N_VDD_XI9.XI106.XI9.MM1_s N_VDD_XI9.XI103.XI1.MM1_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9.XI101.XI9.MM1 N_XI9.XI101.NET43_XI9.XI101.XI9.MM1_d
+ N_ACC3_XI9.XI101.XI9.MM1_g N_VDD_XI9.XI101.XI9.MM1_s N_VDD_XI9.XI102.XI1.MM1_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9.XI86.XI9.MM1 N_XI9.XI86.NET43_XI9.XI86.XI9.MM1_d N_ACC2_XI9.XI86.XI9.MM1_g
+ N_VDD_XI9.XI86.XI9.MM1_s N_VDD_XI9.XI88.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9.XI80.XI9.MM1 N_XI9.XI80.NET43_XI9.XI80.XI9.MM1_d N_ACC1_XI9.XI80.XI9.MM1_g
+ N_VDD_XI9.XI80.XI9.MM1_s N_VDD_XI9.XI82.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9.XI26.XI9.MM1 N_XI9.XI26.NET43_XI9.XI26.XI9.MM1_d N_ACC0_XI9.XI26.XI9.MM1_g
+ N_VDD_XI9.XI26.XI9.MM1_s N_VDD_XI9.XI97.XI4.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9.XI168.XI1.XI1.MM1 N_XI9.XI168.XI1.NET6_XI9.XI168.XI1.XI1.MM1_d
+ N_XI9.NET138_XI9.XI168.XI1.XI1.MM1_g N_VDD_XI9.XI168.XI1.XI1.MM1_s
+ N_VDD_XI9.XI153.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.35e-13
+ PD=7.4e-07 PS=2.48e-06
mXI9.XI167.XI1.XI1.MM1 N_XI9.XI167.XI1.NET6_XI9.XI167.XI1.XI1.MM1_d
+ N_XI9.NET208_XI9.XI167.XI1.XI1.MM1_g N_VDD_XI9.XI167.XI1.XI1.MM1_s
+ N_VDD_XI9.XI154.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.35e-13
+ PD=7.4e-07 PS=2.48e-06
mXI9.XI166.XI1.XI1.MM1 N_XI9.XI166.XI1.NET6_XI9.XI166.XI1.XI1.MM1_d
+ N_XI9.NET202_XI9.XI166.XI1.XI1.MM1_g N_VDD_XI9.XI166.XI1.XI1.MM1_s
+ N_VDD_XI9.XI157.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.35e-13
+ PD=7.4e-07 PS=2.48e-06
mXI9.XI165.XI1.XI1.MM1 N_XI9.XI165.XI1.NET6_XI9.XI165.XI1.XI1.MM1_d
+ N_XI9.NET198_XI9.XI165.XI1.XI1.MM1_g N_VDD_XI9.XI165.XI1.XI1.MM1_s
+ N_VDD_XI9.XI156.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.35e-13
+ PD=7.4e-07 PS=2.48e-06
mXI9.XI159.XI1.XI1.MM1 N_XI9.XI159.XI1.NET6_XI9.XI159.XI1.XI1.MM1_d
+ N_XI9.NET102_XI9.XI159.XI1.XI1.MM1_g N_VDD_XI9.XI159.XI1.XI1.MM1_s
+ N_VDD_XI9.XI155.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.35e-13
+ PD=7.4e-07 PS=2.48e-06
mXI9.XI160.XI1.XI1.MM1 N_XI9.XI160.XI1.NET6_XI9.XI160.XI1.XI1.MM1_d
+ N_XI9.NET108_XI9.XI160.XI1.XI1.MM1_g N_VDD_XI9.XI160.XI1.XI1.MM1_s
+ N_VDD_XI9.XI133.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.35e-13
+ PD=7.4e-07 PS=2.48e-06
mXI9.XI161.XI1.XI1.MM1 N_XI9.XI161.XI1.NET6_XI9.XI161.XI1.XI1.MM1_d
+ N_XI9.NET96_XI9.XI161.XI1.XI1.MM1_g N_VDD_XI9.XI161.XI1.XI1.MM1_s
+ N_VDD_XI9.XI132.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.35e-13
+ PD=7.4e-07 PS=2.48e-06
mXI9.XI162.XI1.XI1.MM1 N_XI9.XI162.XI1.NET6_XI9.XI162.XI1.XI1.MM1_d
+ N_XI9.NET153_XI9.XI162.XI1.XI1.MM1_g N_VDD_XI9.XI162.XI1.XI1.MM1_s
+ N_VDD_XI9.XI131.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.35e-13
+ PD=7.4e-07 PS=2.48e-06
mXI9.XI121.XI1.XI1.MM1 N_XI9.XI121.XI1.NET6_XI9.XI121.XI1.XI1.MM1_d
+ N_XI9.NET54_XI9.XI121.XI1.XI1.MM1_g N_VDD_XI9.XI121.XI1.XI1.MM1_s
+ N_VDD_XI9.XI111.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.35e-13
+ PD=7.4e-07 PS=2.48e-06
mXI9.XI120.XI1.XI1.MM1 N_XI9.XI120.XI1.NET6_XI9.XI120.XI1.XI1.MM1_d
+ N_XI9.NET66_XI9.XI120.XI1.XI1.MM1_g N_VDD_XI9.XI120.XI1.XI1.MM1_s
+ N_VDD_XI9.XI110.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.35e-13
+ PD=7.4e-07 PS=2.48e-06
mXI9.XI119.XI1.XI1.MM1 N_XI9.XI119.XI1.NET6_XI9.XI119.XI1.XI1.MM1_d
+ N_XI9.NET72_XI9.XI119.XI1.XI1.MM1_g N_VDD_XI9.XI119.XI1.XI1.MM1_s
+ N_VDD_XI9.XI103.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.35e-13
+ PD=7.4e-07 PS=2.48e-06
mXI9.XI118.XI1.XI1.MM1 N_XI9.XI118.XI1.NET6_XI9.XI118.XI1.XI1.MM1_d
+ N_XI9.NET60_XI9.XI118.XI1.XI1.MM1_g N_VDD_XI9.XI118.XI1.XI1.MM1_s
+ N_VDD_XI9.XI102.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.35e-13
+ PD=7.4e-07 PS=2.48e-06
mXI9.XI91.XI1.XI1.MM1 N_XI9.XI91.XI1.NET6_XI9.XI91.XI1.XI1.MM1_d
+ N_XI9.NET183_XI9.XI91.XI1.XI1.MM1_g N_VDD_XI9.XI91.XI1.XI1.MM1_s
+ N_VDD_XI9.XI88.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.35e-13
+ PD=7.4e-07 PS=2.48e-06
mXI9.XI90.XI1.XI1.MM1 N_XI9.XI90.XI1.NET6_XI9.XI90.XI1.XI1.MM1_d
+ N_XI9.NET178_XI9.XI90.XI1.XI1.MM1_g N_VDD_XI9.XI90.XI1.XI1.MM1_s
+ N_VDD_XI9.XI82.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.35e-13
+ PD=7.4e-07 PS=2.48e-06
mXI9.XI89.XI1.XI1.MM1 N_XI9.XI89.XI1.NET6_XI9.XI89.XI1.XI1.MM1_d
+ N_CIN1_XI9.XI89.XI1.XI1.MM1_g N_VDD_XI9.XI89.XI1.XI1.MM1_s
+ N_VDD_XI9.XI97.XI4.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.35e-13
+ PD=7.4e-07 PS=2.48e-06
mXI9.XI168.XI1.XI1.MM3 N_XI9.XI168.XI1.NET6_XI9.XI168.XI1.XI1.MM3_d
+ N_XI9.P15_XI9.XI168.XI1.XI1.MM3_g N_VDD_XI9.XI168.XI1.XI1.MM3_s
+ N_VDD_XI9.XI153.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.65e-13
+ PD=7.4e-07 PS=2.52e-06
mXI9.XI167.XI1.XI1.MM3 N_XI9.XI167.XI1.NET6_XI9.XI167.XI1.XI1.MM3_d
+ N_XI9.P14_XI9.XI167.XI1.XI1.MM3_g N_VDD_XI9.XI167.XI1.XI1.MM3_s
+ N_VDD_XI9.XI154.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.65e-13
+ PD=7.4e-07 PS=2.52e-06
mXI9.XI166.XI1.XI1.MM3 N_XI9.XI166.XI1.NET6_XI9.XI166.XI1.XI1.MM3_d
+ N_XI9.P13_XI9.XI166.XI1.XI1.MM3_g N_VDD_XI9.XI166.XI1.XI1.MM3_s
+ N_VDD_XI9.XI157.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.65e-13
+ PD=7.4e-07 PS=2.52e-06
mXI9.XI165.XI1.XI1.MM3 N_XI9.XI165.XI1.NET6_XI9.XI165.XI1.XI1.MM3_d
+ N_XI9.P12_XI9.XI165.XI1.XI1.MM3_g N_VDD_XI9.XI165.XI1.XI1.MM3_s
+ N_VDD_XI9.XI156.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.65e-13
+ PD=7.4e-07 PS=2.52e-06
mXI9.XI159.XI1.XI1.MM3 N_XI9.XI159.XI1.NET6_XI9.XI159.XI1.XI1.MM3_d
+ N_XI9.P11_XI9.XI159.XI1.XI1.MM3_g N_VDD_XI9.XI159.XI1.XI1.MM3_s
+ N_VDD_XI9.XI155.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.65e-13
+ PD=7.4e-07 PS=2.52e-06
mXI9.XI160.XI1.XI1.MM3 N_XI9.XI160.XI1.NET6_XI9.XI160.XI1.XI1.MM3_d
+ N_XI9.P10_XI9.XI160.XI1.XI1.MM3_g N_VDD_XI9.XI160.XI1.XI1.MM3_s
+ N_VDD_XI9.XI133.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.65e-13
+ PD=7.4e-07 PS=2.52e-06
mXI9.XI161.XI1.XI1.MM3 N_XI9.XI161.XI1.NET6_XI9.XI161.XI1.XI1.MM3_d
+ N_XI9.P9_XI9.XI161.XI1.XI1.MM3_g N_VDD_XI9.XI161.XI1.XI1.MM3_s
+ N_VDD_XI9.XI132.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.65e-13
+ PD=7.4e-07 PS=2.52e-06
mXI9.XI162.XI1.XI1.MM3 N_XI9.XI162.XI1.NET6_XI9.XI162.XI1.XI1.MM3_d
+ N_XI9.P8_XI9.XI162.XI1.XI1.MM3_g N_VDD_XI9.XI162.XI1.XI1.MM3_s
+ N_VDD_XI9.XI131.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.65e-13
+ PD=7.4e-07 PS=2.52e-06
mXI9.XI121.XI1.XI1.MM3 N_XI9.XI121.XI1.NET6_XI9.XI121.XI1.XI1.MM3_d
+ N_XI9.P7_XI9.XI121.XI1.XI1.MM3_g N_VDD_XI9.XI121.XI1.XI1.MM3_s
+ N_VDD_XI9.XI111.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.65e-13
+ PD=7.4e-07 PS=2.52e-06
mXI9.XI120.XI1.XI1.MM3 N_XI9.XI120.XI1.NET6_XI9.XI120.XI1.XI1.MM3_d
+ N_XI9.P6_XI9.XI120.XI1.XI1.MM3_g N_VDD_XI9.XI120.XI1.XI1.MM3_s
+ N_VDD_XI9.XI110.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.65e-13
+ PD=7.4e-07 PS=2.52e-06
mXI9.XI119.XI1.XI1.MM3 N_XI9.XI119.XI1.NET6_XI9.XI119.XI1.XI1.MM3_d
+ N_XI9.P5_XI9.XI119.XI1.XI1.MM3_g N_VDD_XI9.XI119.XI1.XI1.MM3_s
+ N_VDD_XI9.XI103.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.65e-13
+ PD=7.4e-07 PS=2.52e-06
mXI9.XI118.XI1.XI1.MM3 N_XI9.XI118.XI1.NET6_XI9.XI118.XI1.XI1.MM3_d
+ N_XI9.P4_XI9.XI118.XI1.XI1.MM3_g N_VDD_XI9.XI118.XI1.XI1.MM3_s
+ N_VDD_XI9.XI102.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.65e-13
+ PD=7.4e-07 PS=2.52e-06
mXI9.XI91.XI1.XI1.MM3 N_XI9.XI91.XI1.NET6_XI9.XI91.XI1.XI1.MM3_d
+ N_XI9.P3_XI9.XI91.XI1.XI1.MM3_g N_VDD_XI9.XI91.XI1.XI1.MM3_s
+ N_VDD_XI9.XI88.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.65e-13
+ PD=7.4e-07 PS=2.52e-06
mXI9.XI90.XI1.XI1.MM3 N_XI9.XI90.XI1.NET6_XI9.XI90.XI1.XI1.MM3_d
+ N_XI9.P2_XI9.XI90.XI1.XI1.MM3_g N_VDD_XI9.XI90.XI1.XI1.MM3_s
+ N_VDD_XI9.XI82.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.65e-13
+ PD=7.4e-07 PS=2.52e-06
mXI9.XI89.XI1.XI1.MM3 N_XI9.XI89.XI1.NET6_XI9.XI89.XI1.XI1.MM3_d
+ N_XI9.P1_XI9.XI89.XI1.XI1.MM3_g N_VDD_XI9.XI89.XI1.XI1.MM3_s
+ N_VDD_XI9.XI97.XI4.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.65e-13
+ PD=7.4e-07 PS=2.52e-06
mXI27.MM1 N_NET214_XI27.MM1_d N_NET218_XI27.MM1_g N_VDD_XI27.MM1_s
+ N_VDD_XI27.MM1_b P_18 L=1.8e-07 W=4.5e-06 AD=2.205e-12 AS=2.205e-12
+ PD=5.48e-06 PS=5.48e-06
mXI28.MM1 N_NET210_XI28.MM1_d N_NET214_XI28.MM1_g N_VDD_XI28.MM1_s
+ N_VDD_XI28.MM1_b P_18 L=1.8e-07 W=9e-06 AD=4.41e-12 AS=4.41e-12 PD=9.98e-06
+ PS=9.98e-06
mXI29.MM1 N_NET222_XI29.MM1_d N_NET210_XI29.MM1_g N_VDD_XI29.MM1_s
+ N_VDD_XI28.MM1_b P_18 L=1.8e-07 W=9e-06 AD=4.41e-12 AS=4.41e-12 PD=9.98e-06
+ PS=9.98e-06
mXI9.XI168.XI1.XI0.MM1 N_XI9.XI168.NET13_XI9.XI168.XI1.XI0.MM1_d
+ N_XI9.XI168.XI1.NET6_XI9.XI168.XI1.XI0.MM1_g N_VDD_XI9.XI168.XI1.XI0.MM1_s
+ N_VDD_XI9.XI153.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI9.XI167.XI1.XI0.MM1 N_XI9.XI167.NET13_XI9.XI167.XI1.XI0.MM1_d
+ N_XI9.XI167.XI1.NET6_XI9.XI167.XI1.XI0.MM1_g N_VDD_XI9.XI167.XI1.XI0.MM1_s
+ N_VDD_XI9.XI154.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI9.XI166.XI1.XI0.MM1 N_XI9.XI166.NET13_XI9.XI166.XI1.XI0.MM1_d
+ N_XI9.XI166.XI1.NET6_XI9.XI166.XI1.XI0.MM1_g N_VDD_XI9.XI166.XI1.XI0.MM1_s
+ N_VDD_XI9.XI157.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI9.XI165.XI1.XI0.MM1 N_XI9.XI165.NET13_XI9.XI165.XI1.XI0.MM1_d
+ N_XI9.XI165.XI1.NET6_XI9.XI165.XI1.XI0.MM1_g N_VDD_XI9.XI165.XI1.XI0.MM1_s
+ N_VDD_XI9.XI156.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI9.XI159.XI1.XI0.MM1 N_XI9.XI159.NET13_XI9.XI159.XI1.XI0.MM1_d
+ N_XI9.XI159.XI1.NET6_XI9.XI159.XI1.XI0.MM1_g N_VDD_XI9.XI159.XI1.XI0.MM1_s
+ N_VDD_XI9.XI155.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI9.XI160.XI1.XI0.MM1 N_XI9.XI160.NET13_XI9.XI160.XI1.XI0.MM1_d
+ N_XI9.XI160.XI1.NET6_XI9.XI160.XI1.XI0.MM1_g N_VDD_XI9.XI160.XI1.XI0.MM1_s
+ N_VDD_XI9.XI133.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI9.XI161.XI1.XI0.MM1 N_XI9.XI161.NET13_XI9.XI161.XI1.XI0.MM1_d
+ N_XI9.XI161.XI1.NET6_XI9.XI161.XI1.XI0.MM1_g N_VDD_XI9.XI161.XI1.XI0.MM1_s
+ N_VDD_XI9.XI132.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI9.XI162.XI1.XI0.MM1 N_XI9.XI162.NET13_XI9.XI162.XI1.XI0.MM1_d
+ N_XI9.XI162.XI1.NET6_XI9.XI162.XI1.XI0.MM1_g N_VDD_XI9.XI162.XI1.XI0.MM1_s
+ N_VDD_XI9.XI131.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI9.XI121.XI1.XI0.MM1 N_XI9.XI121.NET13_XI9.XI121.XI1.XI0.MM1_d
+ N_XI9.XI121.XI1.NET6_XI9.XI121.XI1.XI0.MM1_g N_VDD_XI9.XI121.XI1.XI0.MM1_s
+ N_VDD_XI9.XI111.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI9.XI120.XI1.XI0.MM1 N_XI9.XI120.NET13_XI9.XI120.XI1.XI0.MM1_d
+ N_XI9.XI120.XI1.NET6_XI9.XI120.XI1.XI0.MM1_g N_VDD_XI9.XI120.XI1.XI0.MM1_s
+ N_VDD_XI9.XI110.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI9.XI119.XI1.XI0.MM1 N_XI9.XI119.NET13_XI9.XI119.XI1.XI0.MM1_d
+ N_XI9.XI119.XI1.NET6_XI9.XI119.XI1.XI0.MM1_g N_VDD_XI9.XI119.XI1.XI0.MM1_s
+ N_VDD_XI9.XI103.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI9.XI118.XI1.XI0.MM1 N_XI9.XI118.NET13_XI9.XI118.XI1.XI0.MM1_d
+ N_XI9.XI118.XI1.NET6_XI9.XI118.XI1.XI0.MM1_g N_VDD_XI9.XI118.XI1.XI0.MM1_s
+ N_VDD_XI9.XI102.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI9.XI91.XI1.XI0.MM1 N_XI9.XI91.NET13_XI9.XI91.XI1.XI0.MM1_d
+ N_XI9.XI91.XI1.NET6_XI9.XI91.XI1.XI0.MM1_g N_VDD_XI9.XI91.XI1.XI0.MM1_s
+ N_VDD_XI9.XI88.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI9.XI90.XI1.XI0.MM1 N_XI9.XI90.NET13_XI9.XI90.XI1.XI0.MM1_d
+ N_XI9.XI90.XI1.NET6_XI9.XI90.XI1.XI0.MM1_g N_VDD_XI9.XI90.XI1.XI0.MM1_s
+ N_VDD_XI9.XI82.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI9.XI89.XI1.XI0.MM1 N_XI9.XI89.NET13_XI9.XI89.XI1.XI0.MM1_d
+ N_XI9.XI89.XI1.NET6_XI9.XI89.XI1.XI0.MM1_g N_VDD_XI9.XI89.XI1.XI0.MM1_s
+ N_VDD_XI9.XI97.XI4.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI26.MM1 N_NET218_XI26.MM1_d N_CLK_XI26.MM1_g N_VDD_XI26.MM1_s N_VDD_XI27.MM1_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9.XI168.XI0.XI0.MM1 N_XI9.XI168.XI0.XI0.NET17_XI9.XI168.XI0.XI0.MM1_d
+ N_XI9.XI168.NET13_XI9.XI168.XI0.XI0.MM1_g N_VDD_XI9.XI168.XI0.XI0.MM1_s
+ N_VDD_XI9.XI153.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=4.125e-13 AS=7.35e-13
+ PD=5.5e-07 PS=2.48e-06
mXI9.XI167.XI0.XI0.MM1 N_XI9.XI167.XI0.XI0.NET17_XI9.XI167.XI0.XI0.MM1_d
+ N_XI9.XI167.NET13_XI9.XI167.XI0.XI0.MM1_g N_VDD_XI9.XI167.XI0.XI0.MM1_s
+ N_VDD_XI9.XI154.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=4.125e-13 AS=7.35e-13
+ PD=5.5e-07 PS=2.48e-06
mXI9.XI166.XI0.XI0.MM1 N_XI9.XI166.XI0.XI0.NET17_XI9.XI166.XI0.XI0.MM1_d
+ N_XI9.XI166.NET13_XI9.XI166.XI0.XI0.MM1_g N_VDD_XI9.XI166.XI0.XI0.MM1_s
+ N_VDD_XI9.XI157.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=4.125e-13 AS=7.35e-13
+ PD=5.5e-07 PS=2.48e-06
mXI9.XI165.XI0.XI0.MM1 N_XI9.XI165.XI0.XI0.NET17_XI9.XI165.XI0.XI0.MM1_d
+ N_XI9.XI165.NET13_XI9.XI165.XI0.XI0.MM1_g N_VDD_XI9.XI165.XI0.XI0.MM1_s
+ N_VDD_XI9.XI156.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=4.125e-13 AS=7.35e-13
+ PD=5.5e-07 PS=2.48e-06
mXI9.XI159.XI0.XI0.MM1 N_XI9.XI159.XI0.XI0.NET17_XI9.XI159.XI0.XI0.MM1_d
+ N_XI9.XI159.NET13_XI9.XI159.XI0.XI0.MM1_g N_VDD_XI9.XI159.XI0.XI0.MM1_s
+ N_VDD_XI9.XI155.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=4.125e-13 AS=7.35e-13
+ PD=5.5e-07 PS=2.48e-06
mXI9.XI160.XI0.XI0.MM1 N_XI9.XI160.XI0.XI0.NET17_XI9.XI160.XI0.XI0.MM1_d
+ N_XI9.XI160.NET13_XI9.XI160.XI0.XI0.MM1_g N_VDD_XI9.XI160.XI0.XI0.MM1_s
+ N_VDD_XI9.XI133.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=4.125e-13 AS=7.35e-13
+ PD=5.5e-07 PS=2.48e-06
mXI9.XI161.XI0.XI0.MM1 N_XI9.XI161.XI0.XI0.NET17_XI9.XI161.XI0.XI0.MM1_d
+ N_XI9.XI161.NET13_XI9.XI161.XI0.XI0.MM1_g N_VDD_XI9.XI161.XI0.XI0.MM1_s
+ N_VDD_XI9.XI132.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=4.125e-13 AS=7.35e-13
+ PD=5.5e-07 PS=2.48e-06
mXI9.XI162.XI0.XI0.MM1 N_XI9.XI162.XI0.XI0.NET17_XI9.XI162.XI0.XI0.MM1_d
+ N_XI9.XI162.NET13_XI9.XI162.XI0.XI0.MM1_g N_VDD_XI9.XI162.XI0.XI0.MM1_s
+ N_VDD_XI9.XI131.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=4.125e-13 AS=7.35e-13
+ PD=5.5e-07 PS=2.48e-06
mXI9.XI121.XI0.XI0.MM1 N_XI9.XI121.XI0.XI0.NET17_XI9.XI121.XI0.XI0.MM1_d
+ N_XI9.XI121.NET13_XI9.XI121.XI0.XI0.MM1_g N_VDD_XI9.XI121.XI0.XI0.MM1_s
+ N_VDD_XI9.XI111.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=4.125e-13 AS=7.35e-13
+ PD=5.5e-07 PS=2.48e-06
mXI9.XI120.XI0.XI0.MM1 N_XI9.XI120.XI0.XI0.NET17_XI9.XI120.XI0.XI0.MM1_d
+ N_XI9.XI120.NET13_XI9.XI120.XI0.XI0.MM1_g N_VDD_XI9.XI120.XI0.XI0.MM1_s
+ N_VDD_XI9.XI110.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=4.125e-13 AS=7.35e-13
+ PD=5.5e-07 PS=2.48e-06
mXI9.XI119.XI0.XI0.MM1 N_XI9.XI119.XI0.XI0.NET17_XI9.XI119.XI0.XI0.MM1_d
+ N_XI9.XI119.NET13_XI9.XI119.XI0.XI0.MM1_g N_VDD_XI9.XI119.XI0.XI0.MM1_s
+ N_VDD_XI9.XI103.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=4.125e-13 AS=7.35e-13
+ PD=5.5e-07 PS=2.48e-06
mXI9.XI118.XI0.XI0.MM1 N_XI9.XI118.XI0.XI0.NET17_XI9.XI118.XI0.XI0.MM1_d
+ N_XI9.XI118.NET13_XI9.XI118.XI0.XI0.MM1_g N_VDD_XI9.XI118.XI0.XI0.MM1_s
+ N_VDD_XI9.XI102.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=4.125e-13 AS=7.35e-13
+ PD=5.5e-07 PS=2.48e-06
mXI9.XI91.XI0.XI0.MM1 N_XI9.XI91.XI0.XI0.NET17_XI9.XI91.XI0.XI0.MM1_d
+ N_XI9.XI91.NET13_XI9.XI91.XI0.XI0.MM1_g N_VDD_XI9.XI91.XI0.XI0.MM1_s
+ N_VDD_XI9.XI88.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=4.125e-13 AS=7.35e-13
+ PD=5.5e-07 PS=2.48e-06
mXI9.XI90.XI0.XI0.MM1 N_XI9.XI90.XI0.XI0.NET17_XI9.XI90.XI0.XI0.MM1_d
+ N_XI9.XI90.NET13_XI9.XI90.XI0.XI0.MM1_g N_VDD_XI9.XI90.XI0.XI0.MM1_s
+ N_VDD_XI9.XI82.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=4.125e-13 AS=7.35e-13
+ PD=5.5e-07 PS=2.48e-06
mXI9.XI89.XI0.XI0.MM1 N_XI9.XI89.XI0.XI0.NET17_XI9.XI89.XI0.XI0.MM1_d
+ N_XI9.XI89.NET13_XI9.XI89.XI0.XI0.MM1_g N_VDD_XI9.XI89.XI0.XI0.MM1_s
+ N_VDD_XI9.XI97.XI4.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=4.125e-13 AS=7.35e-13
+ PD=5.5e-07 PS=2.48e-06
mXI9.XI168.XI0.XI0.MM3 N_XI9.XI168.XI0.NET12_XI9.XI168.XI0.XI0.MM3_d
+ N_XI9.G15_XI9.XI168.XI0.XI0.MM3_g
+ N_XI9.XI168.XI0.XI0.NET17_XI9.XI168.XI0.XI0.MM3_s N_VDD_XI9.XI153.XI1.MM1_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=4.125e-13 PD=2.52e-06 PS=5.5e-07
mXI9.XI167.XI0.XI0.MM3 N_XI9.XI167.XI0.NET12_XI9.XI167.XI0.XI0.MM3_d
+ N_XI9.G14_XI9.XI167.XI0.XI0.MM3_g
+ N_XI9.XI167.XI0.XI0.NET17_XI9.XI167.XI0.XI0.MM3_s N_VDD_XI9.XI154.XI1.MM1_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=4.125e-13 PD=2.52e-06 PS=5.5e-07
mXI9.XI166.XI0.XI0.MM3 N_XI9.XI166.XI0.NET12_XI9.XI166.XI0.XI0.MM3_d
+ N_XI9.G13_XI9.XI166.XI0.XI0.MM3_g
+ N_XI9.XI166.XI0.XI0.NET17_XI9.XI166.XI0.XI0.MM3_s N_VDD_XI9.XI157.XI1.MM1_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=4.125e-13 PD=2.52e-06 PS=5.5e-07
mXI9.XI165.XI0.XI0.MM3 N_XI9.XI165.XI0.NET12_XI9.XI165.XI0.XI0.MM3_d
+ N_XI9.G12_XI9.XI165.XI0.XI0.MM3_g
+ N_XI9.XI165.XI0.XI0.NET17_XI9.XI165.XI0.XI0.MM3_s N_VDD_XI9.XI156.XI1.MM1_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=4.125e-13 PD=2.52e-06 PS=5.5e-07
mXI9.XI159.XI0.XI0.MM3 N_XI9.XI159.XI0.NET12_XI9.XI159.XI0.XI0.MM3_d
+ N_XI9.G11_XI9.XI159.XI0.XI0.MM3_g
+ N_XI9.XI159.XI0.XI0.NET17_XI9.XI159.XI0.XI0.MM3_s N_VDD_XI9.XI155.XI1.MM1_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=4.125e-13 PD=2.52e-06 PS=5.5e-07
mXI9.XI160.XI0.XI0.MM3 N_XI9.XI160.XI0.NET12_XI9.XI160.XI0.XI0.MM3_d
+ N_XI9.G10_XI9.XI160.XI0.XI0.MM3_g
+ N_XI9.XI160.XI0.XI0.NET17_XI9.XI160.XI0.XI0.MM3_s N_VDD_XI9.XI133.XI1.MM1_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=4.125e-13 PD=2.52e-06 PS=5.5e-07
mXI9.XI161.XI0.XI0.MM3 N_XI9.XI161.XI0.NET12_XI9.XI161.XI0.XI0.MM3_d
+ N_XI9.G9_XI9.XI161.XI0.XI0.MM3_g
+ N_XI9.XI161.XI0.XI0.NET17_XI9.XI161.XI0.XI0.MM3_s N_VDD_XI9.XI132.XI1.MM1_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=4.125e-13 PD=2.52e-06 PS=5.5e-07
mXI9.XI162.XI0.XI0.MM3 N_XI9.XI162.XI0.NET12_XI9.XI162.XI0.XI0.MM3_d
+ N_XI9.G8_XI9.XI162.XI0.XI0.MM3_g
+ N_XI9.XI162.XI0.XI0.NET17_XI9.XI162.XI0.XI0.MM3_s N_VDD_XI9.XI131.XI1.MM1_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=4.125e-13 PD=2.52e-06 PS=5.5e-07
mXI9.XI121.XI0.XI0.MM3 N_XI9.XI121.XI0.NET12_XI9.XI121.XI0.XI0.MM3_d
+ N_XI9.G7_XI9.XI121.XI0.XI0.MM3_g
+ N_XI9.XI121.XI0.XI0.NET17_XI9.XI121.XI0.XI0.MM3_s N_VDD_XI9.XI111.XI1.MM1_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=4.125e-13 PD=2.52e-06 PS=5.5e-07
mXI9.XI120.XI0.XI0.MM3 N_XI9.XI120.XI0.NET12_XI9.XI120.XI0.XI0.MM3_d
+ N_XI9.G6_XI9.XI120.XI0.XI0.MM3_g
+ N_XI9.XI120.XI0.XI0.NET17_XI9.XI120.XI0.XI0.MM3_s N_VDD_XI9.XI110.XI1.MM1_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=4.125e-13 PD=2.52e-06 PS=5.5e-07
mXI9.XI119.XI0.XI0.MM3 N_XI9.XI119.XI0.NET12_XI9.XI119.XI0.XI0.MM3_d
+ N_XI9.G5_XI9.XI119.XI0.XI0.MM3_g
+ N_XI9.XI119.XI0.XI0.NET17_XI9.XI119.XI0.XI0.MM3_s N_VDD_XI9.XI103.XI1.MM1_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=4.125e-13 PD=2.52e-06 PS=5.5e-07
mXI9.XI118.XI0.XI0.MM3 N_XI9.XI118.XI0.NET12_XI9.XI118.XI0.XI0.MM3_d
+ N_XI9.G4_XI9.XI118.XI0.XI0.MM3_g
+ N_XI9.XI118.XI0.XI0.NET17_XI9.XI118.XI0.XI0.MM3_s N_VDD_XI9.XI102.XI1.MM1_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=4.125e-13 PD=2.52e-06 PS=5.5e-07
mXI9.XI91.XI0.XI0.MM3 N_XI9.XI91.XI0.NET12_XI9.XI91.XI0.XI0.MM3_d
+ N_XI9.G3_XI9.XI91.XI0.XI0.MM3_g
+ N_XI9.XI91.XI0.XI0.NET17_XI9.XI91.XI0.XI0.MM3_s N_VDD_XI9.XI88.XI1.MM1_b P_18
+ L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=4.125e-13 PD=2.52e-06 PS=5.5e-07
mXI9.XI90.XI0.XI0.MM3 N_XI9.XI90.XI0.NET12_XI9.XI90.XI0.XI0.MM3_d
+ N_XI9.G2_XI9.XI90.XI0.XI0.MM3_g
+ N_XI9.XI90.XI0.XI0.NET17_XI9.XI90.XI0.XI0.MM3_s N_VDD_XI9.XI82.XI1.MM1_b P_18
+ L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=4.125e-13 PD=2.52e-06 PS=5.5e-07
mXI9.XI89.XI0.XI0.MM3 N_XI9.XI89.XI0.NET12_XI9.XI89.XI0.XI0.MM3_d
+ N_XI9.G1_XI9.XI89.XI0.XI0.MM3_g
+ N_XI9.XI89.XI0.XI0.NET17_XI9.XI89.XI0.XI0.MM3_s N_VDD_XI9.XI97.XI4.MM1_b P_18
+ L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=4.125e-13 PD=2.52e-06 PS=5.5e-07
mXI9.XI168.XI0.XI1.MM1 N_XI9.NET298_XI9.XI168.XI0.XI1.MM1_d
+ N_XI9.XI168.XI0.NET12_XI9.XI168.XI0.XI1.MM1_g N_VDD_XI9.XI168.XI0.XI1.MM1_s
+ N_VDD_XI9.XI153.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI9.XI167.XI0.XI1.MM1 N_XI9.NET138_XI9.XI167.XI0.XI1.MM1_d
+ N_XI9.XI167.XI0.NET12_XI9.XI167.XI0.XI1.MM1_g N_VDD_XI9.XI167.XI0.XI1.MM1_s
+ N_VDD_XI9.XI154.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI9.XI166.XI0.XI1.MM1 N_XI9.NET208_XI9.XI166.XI0.XI1.MM1_d
+ N_XI9.XI166.XI0.NET12_XI9.XI166.XI0.XI1.MM1_g N_VDD_XI9.XI166.XI0.XI1.MM1_s
+ N_VDD_XI9.XI157.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI9.XI165.XI0.XI1.MM1 N_XI9.NET202_XI9.XI165.XI0.XI1.MM1_d
+ N_XI9.XI165.XI0.NET12_XI9.XI165.XI0.XI1.MM1_g N_VDD_XI9.XI165.XI0.XI1.MM1_s
+ N_VDD_XI9.XI156.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI9.XI159.XI0.XI1.MM1 N_XI9.NET198_XI9.XI159.XI0.XI1.MM1_d
+ N_XI9.XI159.XI0.NET12_XI9.XI159.XI0.XI1.MM1_g N_VDD_XI9.XI159.XI0.XI1.MM1_s
+ N_VDD_XI9.XI155.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI9.XI160.XI0.XI1.MM1 N_XI9.NET102_XI9.XI160.XI0.XI1.MM1_d
+ N_XI9.XI160.XI0.NET12_XI9.XI160.XI0.XI1.MM1_g N_VDD_XI9.XI160.XI0.XI1.MM1_s
+ N_VDD_XI9.XI133.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI9.XI161.XI0.XI1.MM1 N_XI9.NET108_XI9.XI161.XI0.XI1.MM1_d
+ N_XI9.XI161.XI0.NET12_XI9.XI161.XI0.XI1.MM1_g N_VDD_XI9.XI161.XI0.XI1.MM1_s
+ N_VDD_XI9.XI132.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI9.XI162.XI0.XI1.MM1 N_XI9.NET96_XI9.XI162.XI0.XI1.MM1_d
+ N_XI9.XI162.XI0.NET12_XI9.XI162.XI0.XI1.MM1_g N_VDD_XI9.XI162.XI0.XI1.MM1_s
+ N_VDD_XI9.XI131.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI9.XI121.XI0.XI1.MM1 N_XI9.NET153_XI9.XI121.XI0.XI1.MM1_d
+ N_XI9.XI121.XI0.NET12_XI9.XI121.XI0.XI1.MM1_g N_VDD_XI9.XI121.XI0.XI1.MM1_s
+ N_VDD_XI9.XI111.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI9.XI120.XI0.XI1.MM1 N_XI9.NET54_XI9.XI120.XI0.XI1.MM1_d
+ N_XI9.XI120.XI0.NET12_XI9.XI120.XI0.XI1.MM1_g N_VDD_XI9.XI120.XI0.XI1.MM1_s
+ N_VDD_XI9.XI110.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI9.XI119.XI0.XI1.MM1 N_XI9.NET66_XI9.XI119.XI0.XI1.MM1_d
+ N_XI9.XI119.XI0.NET12_XI9.XI119.XI0.XI1.MM1_g N_VDD_XI9.XI119.XI0.XI1.MM1_s
+ N_VDD_XI9.XI103.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI9.XI118.XI0.XI1.MM1 N_XI9.NET72_XI9.XI118.XI0.XI1.MM1_d
+ N_XI9.XI118.XI0.NET12_XI9.XI118.XI0.XI1.MM1_g N_VDD_XI9.XI118.XI0.XI1.MM1_s
+ N_VDD_XI9.XI102.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI9.XI91.XI0.XI1.MM1 N_XI9.NET60_XI9.XI91.XI0.XI1.MM1_d
+ N_XI9.XI91.XI0.NET12_XI9.XI91.XI0.XI1.MM1_g N_VDD_XI9.XI91.XI0.XI1.MM1_s
+ N_VDD_XI9.XI88.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI9.XI90.XI0.XI1.MM1 N_XI9.NET183_XI9.XI90.XI0.XI1.MM1_d
+ N_XI9.XI90.XI0.NET12_XI9.XI90.XI0.XI1.MM1_g N_VDD_XI9.XI90.XI0.XI1.MM1_s
+ N_VDD_XI9.XI82.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI9.XI89.XI0.XI1.MM1 N_XI9.NET178_XI9.XI89.XI0.XI1.MM1_d
+ N_XI9.XI89.XI0.NET12_XI9.XI89.XI0.XI1.MM1_g N_VDD_XI9.XI89.XI0.XI1.MM1_s
+ N_VDD_XI9.XI97.XI4.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI9.XI182.XI4.MM1 N_XI9.XI182.NET39_XI9.XI182.XI4.MM1_d
+ N_XI9.NET298_XI9.XI182.XI4.MM1_g N_VDD_XI9.XI182.XI4.MM1_s
+ N_VDD_XI9.XI153.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI9.XI181.XI4.MM1 N_XI9.XI181.NET39_XI9.XI181.XI4.MM1_d
+ N_XI9.NET138_XI9.XI181.XI4.MM1_g N_VDD_XI9.XI181.XI4.MM1_s
+ N_VDD_XI9.XI154.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI9.XI180.XI4.MM1 N_XI9.XI180.NET39_XI9.XI180.XI4.MM1_d
+ N_XI9.NET208_XI9.XI180.XI4.MM1_g N_VDD_XI9.XI180.XI4.MM1_s
+ N_VDD_XI9.XI157.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI9.XI179.XI9.MM1 N_XI9.XI179.NET43_XI9.XI179.XI9.MM1_d
+ N_XI9.NET202_XI9.XI179.XI9.MM1_g N_VDD_XI9.XI179.XI9.MM1_s
+ N_VDD_XI9.XI156.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI9.XI178.XI4.MM1 N_XI9.XI178.NET39_XI9.XI178.XI4.MM1_d
+ N_XI9.NET198_XI9.XI178.XI4.MM1_g N_VDD_XI9.XI178.XI4.MM1_s
+ N_VDD_XI9.XI155.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI9.XI177.XI4.MM1 N_XI9.XI177.NET39_XI9.XI177.XI4.MM1_d
+ N_XI9.NET102_XI9.XI177.XI4.MM1_g N_VDD_XI9.XI177.XI4.MM1_s
+ N_VDD_XI9.XI133.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI9.XI176.XI4.MM1 N_XI9.XI176.NET39_XI9.XI176.XI4.MM1_d
+ N_XI9.NET108_XI9.XI176.XI4.MM1_g N_VDD_XI9.XI176.XI4.MM1_s
+ N_VDD_XI9.XI132.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI9.XI175.XI4.MM1 N_XI9.XI175.NET39_XI9.XI175.XI4.MM1_d
+ N_XI9.NET96_XI9.XI175.XI4.MM1_g N_VDD_XI9.XI175.XI4.MM1_s
+ N_VDD_XI9.XI131.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI9.XI174.XI4.MM1 N_XI9.XI174.NET39_XI9.XI174.XI4.MM1_d
+ N_XI9.NET153_XI9.XI174.XI4.MM1_g N_VDD_XI9.XI174.XI4.MM1_s
+ N_VDD_XI9.XI111.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI9.XI173.XI4.MM1 N_XI9.XI173.NET39_XI9.XI173.XI4.MM1_d
+ N_XI9.NET54_XI9.XI173.XI4.MM1_g N_VDD_XI9.XI173.XI4.MM1_s
+ N_VDD_XI9.XI110.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI9.XI172.XI4.MM1 N_XI9.XI172.NET39_XI9.XI172.XI4.MM1_d
+ N_XI9.NET66_XI9.XI172.XI4.MM1_g N_VDD_XI9.XI172.XI4.MM1_s
+ N_VDD_XI9.XI103.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI9.XI171.XI4.MM1 N_XI9.XI171.NET39_XI9.XI171.XI4.MM1_d
+ N_XI9.NET72_XI9.XI171.XI4.MM1_g N_VDD_XI9.XI171.XI4.MM1_s
+ N_VDD_XI9.XI102.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI9.XI170.XI4.MM1 N_XI9.XI170.NET39_XI9.XI170.XI4.MM1_d
+ N_XI9.NET60_XI9.XI170.XI4.MM1_g N_VDD_XI9.XI170.XI4.MM1_s
+ N_VDD_XI9.XI88.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI9.XI96.XI4.MM1 N_XI9.XI96.NET39_XI9.XI96.XI4.MM1_d
+ N_XI9.NET183_XI9.XI96.XI4.MM1_g N_VDD_XI9.XI96.XI4.MM1_s
+ N_VDD_XI9.XI82.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI9.XI93.XI4.MM1 N_XI9.XI93.NET39_XI9.XI93.XI4.MM1_d
+ N_XI9.NET178_XI9.XI93.XI4.MM1_g N_VDD_XI9.XI93.XI4.MM1_s
+ N_VDD_XI9.XI97.XI4.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI9.XI182.MM3 N_XI9.XI182.NET37_XI9.XI182.MM3_d
+ N_XI9.XI182.NET39_XI9.XI182.MM3_g N_VDD_XI9.XI182.MM3_s
+ N_VDD_XI9.XI153.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=6.7125e-13 AS=9.675e-13
+ PD=8.95e-07 PS=2.79e-06
mXI9.XI181.MM3 N_XI9.XI181.NET37_XI9.XI181.MM3_d
+ N_XI9.XI181.NET39_XI9.XI181.MM3_g N_VDD_XI9.XI181.MM3_s
+ N_VDD_XI9.XI154.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=6.7125e-13 AS=9.675e-13
+ PD=8.95e-07 PS=2.79e-06
mXI9.XI180.MM3 N_XI9.XI180.NET37_XI9.XI180.MM3_d
+ N_XI9.XI180.NET39_XI9.XI180.MM3_g N_VDD_XI9.XI180.MM3_s
+ N_VDD_XI9.XI157.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=6.7125e-13 AS=9.675e-13
+ PD=8.95e-07 PS=2.79e-06
mXI9.XI179.MM5 N_XI9.XI179.NET25_XI9.XI179.MM5_d
+ N_XI9.XI179.NET43_XI9.XI179.MM5_g N_VDD_XI9.XI179.MM5_s
+ N_VDD_XI9.XI156.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=6.7125e-13 AS=9.675e-13
+ PD=8.95e-07 PS=2.79e-06
mXI9.XI178.MM3 N_XI9.XI178.NET37_XI9.XI178.MM3_d
+ N_XI9.XI178.NET39_XI9.XI178.MM3_g N_VDD_XI9.XI178.MM3_s
+ N_VDD_XI9.XI155.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=6.7125e-13 AS=9.675e-13
+ PD=8.95e-07 PS=2.79e-06
mXI9.XI177.MM3 N_XI9.XI177.NET37_XI9.XI177.MM3_d
+ N_XI9.XI177.NET39_XI9.XI177.MM3_g N_VDD_XI9.XI177.MM3_s
+ N_VDD_XI9.XI133.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=6.7125e-13 AS=9.675e-13
+ PD=8.95e-07 PS=2.79e-06
mXI9.XI176.MM3 N_XI9.XI176.NET37_XI9.XI176.MM3_d
+ N_XI9.XI176.NET39_XI9.XI176.MM3_g N_VDD_XI9.XI176.MM3_s
+ N_VDD_XI9.XI132.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=6.7125e-13 AS=9.675e-13
+ PD=8.95e-07 PS=2.79e-06
mXI9.XI175.MM3 N_XI9.XI175.NET37_XI9.XI175.MM3_d
+ N_XI9.XI175.NET39_XI9.XI175.MM3_g N_VDD_XI9.XI175.MM3_s
+ N_VDD_XI9.XI131.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=6.7125e-13 AS=9.675e-13
+ PD=8.95e-07 PS=2.79e-06
mXI9.XI174.MM3 N_XI9.XI174.NET37_XI9.XI174.MM3_d
+ N_XI9.XI174.NET39_XI9.XI174.MM3_g N_VDD_XI9.XI174.MM3_s
+ N_VDD_XI9.XI111.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=6.7125e-13 AS=9.675e-13
+ PD=8.95e-07 PS=2.79e-06
mXI9.XI173.MM3 N_XI9.XI173.NET37_XI9.XI173.MM3_d
+ N_XI9.XI173.NET39_XI9.XI173.MM3_g N_VDD_XI9.XI173.MM3_s
+ N_VDD_XI9.XI110.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=6.7125e-13 AS=9.675e-13
+ PD=8.95e-07 PS=2.79e-06
mXI9.XI172.MM3 N_XI9.XI172.NET37_XI9.XI172.MM3_d
+ N_XI9.XI172.NET39_XI9.XI172.MM3_g N_VDD_XI9.XI172.MM3_s
+ N_VDD_XI9.XI103.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=6.7125e-13 AS=9.675e-13
+ PD=8.95e-07 PS=2.79e-06
mXI9.XI171.MM3 N_XI9.XI171.NET37_XI9.XI171.MM3_d
+ N_XI9.XI171.NET39_XI9.XI171.MM3_g N_VDD_XI9.XI171.MM3_s
+ N_VDD_XI9.XI102.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=6.7125e-13 AS=9.675e-13
+ PD=8.95e-07 PS=2.79e-06
mXI9.XI170.MM3 N_XI9.XI170.NET37_XI9.XI170.MM3_d
+ N_XI9.XI170.NET39_XI9.XI170.MM3_g N_VDD_XI9.XI170.MM3_s
+ N_VDD_XI9.XI88.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=6.7125e-13 AS=9.675e-13
+ PD=8.95e-07 PS=2.79e-06
mXI9.XI96.MM3 N_XI9.XI96.NET37_XI9.XI96.MM3_d N_XI9.XI96.NET39_XI9.XI96.MM3_g
+ N_VDD_XI9.XI96.MM3_s N_VDD_XI9.XI82.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=6.7125e-13 AS=9.675e-13 PD=8.95e-07 PS=2.79e-06
mXI9.XI93.MM3 N_XI9.XI93.NET37_XI9.XI93.MM3_d N_XI9.XI93.NET39_XI9.XI93.MM3_g
+ N_VDD_XI9.XI93.MM3_s N_VDD_XI9.XI97.XI4.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=6.7125e-13 AS=9.675e-13 PD=8.95e-07 PS=2.79e-06
mXI9.XI182.MM1 N_NET177_XI9.XI182.MM1_d N_XI9.P16_XI9.XI182.MM1_g
+ N_XI9.XI182.NET37_XI9.XI182.MM1_s N_VDD_XI9.XI153.XI1.MM1_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.425e-12 AS=6.7125e-13 PD=1.9e-06 PS=8.95e-07
mXI9.XI181.MM1 N_NET178_XI9.XI181.MM1_d N_XI9.P15_XI9.XI181.MM1_g
+ N_XI9.XI181.NET37_XI9.XI181.MM1_s N_VDD_XI9.XI154.XI1.MM1_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.425e-12 AS=6.7125e-13 PD=1.9e-06 PS=8.95e-07
mXI9.XI180.MM1 N_NET179_XI9.XI180.MM1_d N_XI9.P14_XI9.XI180.MM1_g
+ N_XI9.XI180.NET37_XI9.XI180.MM1_s N_VDD_XI9.XI157.XI1.MM1_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.425e-12 AS=6.7125e-13 PD=1.9e-06 PS=8.95e-07
mXI9.XI179.MM4 N_NET180_XI9.XI179.MM4_d N_XI9.P13_XI9.XI179.MM4_g
+ N_XI9.XI179.NET25_XI9.XI179.MM4_s N_VDD_XI9.XI156.XI1.MM1_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.425e-12 AS=6.7125e-13 PD=1.9e-06 PS=8.95e-07
mXI9.XI178.MM1 N_NET181_XI9.XI178.MM1_d N_XI9.P12_XI9.XI178.MM1_g
+ N_XI9.XI178.NET37_XI9.XI178.MM1_s N_VDD_XI9.XI155.XI1.MM1_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.425e-12 AS=6.7125e-13 PD=1.9e-06 PS=8.95e-07
mXI9.XI177.MM1 N_NET182_XI9.XI177.MM1_d N_XI9.P11_XI9.XI177.MM1_g
+ N_XI9.XI177.NET37_XI9.XI177.MM1_s N_VDD_XI9.XI133.XI1.MM1_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.425e-12 AS=6.7125e-13 PD=1.9e-06 PS=8.95e-07
mXI9.XI176.MM1 N_NET183_XI9.XI176.MM1_d N_XI9.P10_XI9.XI176.MM1_g
+ N_XI9.XI176.NET37_XI9.XI176.MM1_s N_VDD_XI9.XI132.XI1.MM1_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.425e-12 AS=6.7125e-13 PD=1.9e-06 PS=8.95e-07
mXI9.XI175.MM1 N_NET184_XI9.XI175.MM1_d N_XI9.P9_XI9.XI175.MM1_g
+ N_XI9.XI175.NET37_XI9.XI175.MM1_s N_VDD_XI9.XI131.XI1.MM1_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.425e-12 AS=6.7125e-13 PD=1.9e-06 PS=8.95e-07
mXI9.XI174.MM1 N_NET185_XI9.XI174.MM1_d N_XI9.P8_XI9.XI174.MM1_g
+ N_XI9.XI174.NET37_XI9.XI174.MM1_s N_VDD_XI9.XI111.XI1.MM1_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.425e-12 AS=6.7125e-13 PD=1.9e-06 PS=8.95e-07
mXI9.XI173.MM1 N_NET186_XI9.XI173.MM1_d N_XI9.P7_XI9.XI173.MM1_g
+ N_XI9.XI173.NET37_XI9.XI173.MM1_s N_VDD_XI9.XI110.XI1.MM1_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.425e-12 AS=6.7125e-13 PD=1.9e-06 PS=8.95e-07
mXI9.XI172.MM1 N_NET187_XI9.XI172.MM1_d N_XI9.P6_XI9.XI172.MM1_g
+ N_XI9.XI172.NET37_XI9.XI172.MM1_s N_VDD_XI9.XI103.XI1.MM1_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.425e-12 AS=6.7125e-13 PD=1.9e-06 PS=8.95e-07
mXI9.XI171.MM1 N_NET188_XI9.XI171.MM1_d N_XI9.P5_XI9.XI171.MM1_g
+ N_XI9.XI171.NET37_XI9.XI171.MM1_s N_VDD_XI9.XI102.XI1.MM1_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.425e-12 AS=6.7125e-13 PD=1.9e-06 PS=8.95e-07
mXI9.XI170.MM1 N_NET189_XI9.XI170.MM1_d N_XI9.P4_XI9.XI170.MM1_g
+ N_XI9.XI170.NET37_XI9.XI170.MM1_s N_VDD_XI9.XI88.XI1.MM1_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.425e-12 AS=6.7125e-13 PD=1.9e-06 PS=8.95e-07
mXI9.XI96.MM1 N_NET190_XI9.XI96.MM1_d N_XI9.P3_XI9.XI96.MM1_g
+ N_XI9.XI96.NET37_XI9.XI96.MM1_s N_VDD_XI9.XI82.XI1.MM1_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.425e-12 AS=6.7125e-13 PD=1.9e-06 PS=8.95e-07
mXI9.XI93.MM1 N_NET191_XI9.XI93.MM1_d N_XI9.P2_XI9.XI93.MM1_g
+ N_XI9.XI93.NET37_XI9.XI93.MM1_s N_VDD_XI9.XI97.XI4.MM1_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.425e-12 AS=6.7125e-13 PD=1.9e-06 PS=8.95e-07
mXI9.XI182.MM5 N_NET177_XI9.XI182.MM5_d N_XI9.XI182.NET43_XI9.XI182.MM5_g
+ N_XI9.XI182.NET25_XI9.XI182.MM5_s N_VDD_XI9.XI153.XI1.MM1_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.425e-12 AS=5.4375e-13 PD=1.9e-06 PS=7.25e-07
mXI9.XI181.MM5 N_NET178_XI9.XI181.MM5_d N_XI9.XI181.NET43_XI9.XI181.MM5_g
+ N_XI9.XI181.NET25_XI9.XI181.MM5_s N_VDD_XI9.XI154.XI1.MM1_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.425e-12 AS=5.4375e-13 PD=1.9e-06 PS=7.25e-07
mXI9.XI180.MM5 N_NET179_XI9.XI180.MM5_d N_XI9.XI180.NET43_XI9.XI180.MM5_g
+ N_XI9.XI180.NET25_XI9.XI180.MM5_s N_VDD_XI9.XI157.XI1.MM1_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.425e-12 AS=5.4375e-13 PD=1.9e-06 PS=7.25e-07
mXI9.XI179.MM3 N_NET180_XI9.XI179.MM3_d N_XI9.XI179.NET39_XI9.XI179.MM3_g
+ N_XI9.XI179.NET37_XI9.XI179.MM3_s N_VDD_XI9.XI156.XI1.MM1_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.425e-12 AS=5.4375e-13 PD=1.9e-06 PS=7.25e-07
mXI9.XI178.MM5 N_NET181_XI9.XI178.MM5_d N_XI9.XI178.NET43_XI9.XI178.MM5_g
+ N_XI9.XI178.NET25_XI9.XI178.MM5_s N_VDD_XI9.XI155.XI1.MM1_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.425e-12 AS=5.4375e-13 PD=1.9e-06 PS=7.25e-07
mXI9.XI177.MM5 N_NET182_XI9.XI177.MM5_d N_XI9.XI177.NET43_XI9.XI177.MM5_g
+ N_XI9.XI177.NET25_XI9.XI177.MM5_s N_VDD_XI9.XI133.XI1.MM1_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.425e-12 AS=5.4375e-13 PD=1.9e-06 PS=7.25e-07
mXI9.XI176.MM5 N_NET183_XI9.XI176.MM5_d N_XI9.XI176.NET43_XI9.XI176.MM5_g
+ N_XI9.XI176.NET25_XI9.XI176.MM5_s N_VDD_XI9.XI132.XI1.MM1_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.425e-12 AS=5.4375e-13 PD=1.9e-06 PS=7.25e-07
mXI9.XI175.MM5 N_NET184_XI9.XI175.MM5_d N_XI9.XI175.NET43_XI9.XI175.MM5_g
+ N_XI9.XI175.NET25_XI9.XI175.MM5_s N_VDD_XI9.XI131.XI1.MM1_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.425e-12 AS=5.4375e-13 PD=1.9e-06 PS=7.25e-07
mXI9.XI174.MM5 N_NET185_XI9.XI174.MM5_d N_XI9.XI174.NET43_XI9.XI174.MM5_g
+ N_XI9.XI174.NET25_XI9.XI174.MM5_s N_VDD_XI9.XI111.XI1.MM1_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.425e-12 AS=5.4375e-13 PD=1.9e-06 PS=7.25e-07
mXI9.XI173.MM5 N_NET186_XI9.XI173.MM5_d N_XI9.XI173.NET43_XI9.XI173.MM5_g
+ N_XI9.XI173.NET25_XI9.XI173.MM5_s N_VDD_XI9.XI110.XI1.MM1_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.425e-12 AS=5.4375e-13 PD=1.9e-06 PS=7.25e-07
mXI9.XI172.MM5 N_NET187_XI9.XI172.MM5_d N_XI9.XI172.NET43_XI9.XI172.MM5_g
+ N_XI9.XI172.NET25_XI9.XI172.MM5_s N_VDD_XI9.XI103.XI1.MM1_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.425e-12 AS=5.4375e-13 PD=1.9e-06 PS=7.25e-07
mXI9.XI171.MM5 N_NET188_XI9.XI171.MM5_d N_XI9.XI171.NET43_XI9.XI171.MM5_g
+ N_XI9.XI171.NET25_XI9.XI171.MM5_s N_VDD_XI9.XI102.XI1.MM1_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.425e-12 AS=5.4375e-13 PD=1.9e-06 PS=7.25e-07
mXI9.XI170.MM5 N_NET189_XI9.XI170.MM5_d N_XI9.XI170.NET43_XI9.XI170.MM5_g
+ N_XI9.XI170.NET25_XI9.XI170.MM5_s N_VDD_XI9.XI88.XI1.MM1_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.425e-12 AS=5.4375e-13 PD=1.9e-06 PS=7.25e-07
mXI9.XI96.MM5 N_NET190_XI9.XI96.MM5_d N_XI9.XI96.NET43_XI9.XI96.MM5_g
+ N_XI9.XI96.NET25_XI9.XI96.MM5_s N_VDD_XI9.XI82.XI1.MM1_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.425e-12 AS=5.4375e-13 PD=1.9e-06 PS=7.25e-07
mXI9.XI93.MM5 N_NET191_XI9.XI93.MM5_d N_XI9.XI93.NET43_XI9.XI93.MM5_g
+ N_XI9.XI93.NET25_XI9.XI93.MM5_s N_VDD_XI9.XI97.XI4.MM1_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.425e-12 AS=5.4375e-13 PD=1.9e-06 PS=7.25e-07
mXI9.XI182.MM4 N_XI9.XI182.NET25_XI9.XI182.MM4_d N_XI9.NET298_XI9.XI182.MM4_g
+ N_VDD_XI9.XI182.MM4_s N_VDD_XI9.XI153.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=5.4375e-13 AS=7.65e-13 PD=7.25e-07 PS=2.52e-06
mXI9.XI181.MM4 N_XI9.XI181.NET25_XI9.XI181.MM4_d N_XI9.NET138_XI9.XI181.MM4_g
+ N_VDD_XI9.XI181.MM4_s N_VDD_XI9.XI154.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=5.4375e-13 AS=7.65e-13 PD=7.25e-07 PS=2.52e-06
mXI9.XI180.MM4 N_XI9.XI180.NET25_XI9.XI180.MM4_d N_XI9.NET208_XI9.XI180.MM4_g
+ N_VDD_XI9.XI180.MM4_s N_VDD_XI9.XI157.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=5.4375e-13 AS=7.65e-13 PD=7.25e-07 PS=2.52e-06
mXI9.XI179.MM1 N_XI9.XI179.NET37_XI9.XI179.MM1_d N_XI9.NET202_XI9.XI179.MM1_g
+ N_VDD_XI9.XI179.MM1_s N_VDD_XI9.XI156.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=5.4375e-13 AS=7.65e-13 PD=7.25e-07 PS=2.52e-06
mXI9.XI178.MM4 N_XI9.XI178.NET25_XI9.XI178.MM4_d N_XI9.NET198_XI9.XI178.MM4_g
+ N_VDD_XI9.XI178.MM4_s N_VDD_XI9.XI155.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=5.4375e-13 AS=7.65e-13 PD=7.25e-07 PS=2.52e-06
mXI9.XI177.MM4 N_XI9.XI177.NET25_XI9.XI177.MM4_d N_XI9.NET102_XI9.XI177.MM4_g
+ N_VDD_XI9.XI177.MM4_s N_VDD_XI9.XI133.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=5.4375e-13 AS=7.65e-13 PD=7.25e-07 PS=2.52e-06
mXI9.XI176.MM4 N_XI9.XI176.NET25_XI9.XI176.MM4_d N_XI9.NET108_XI9.XI176.MM4_g
+ N_VDD_XI9.XI176.MM4_s N_VDD_XI9.XI132.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=5.4375e-13 AS=7.65e-13 PD=7.25e-07 PS=2.52e-06
mXI9.XI175.MM4 N_XI9.XI175.NET25_XI9.XI175.MM4_d N_XI9.NET96_XI9.XI175.MM4_g
+ N_VDD_XI9.XI175.MM4_s N_VDD_XI9.XI131.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=5.4375e-13 AS=7.65e-13 PD=7.25e-07 PS=2.52e-06
mXI9.XI174.MM4 N_XI9.XI174.NET25_XI9.XI174.MM4_d N_XI9.NET153_XI9.XI174.MM4_g
+ N_VDD_XI9.XI174.MM4_s N_VDD_XI9.XI111.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=5.4375e-13 AS=7.65e-13 PD=7.25e-07 PS=2.52e-06
mXI9.XI173.MM4 N_XI9.XI173.NET25_XI9.XI173.MM4_d N_XI9.NET54_XI9.XI173.MM4_g
+ N_VDD_XI9.XI173.MM4_s N_VDD_XI9.XI110.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=5.4375e-13 AS=7.65e-13 PD=7.25e-07 PS=2.52e-06
mXI9.XI172.MM4 N_XI9.XI172.NET25_XI9.XI172.MM4_d N_XI9.NET66_XI9.XI172.MM4_g
+ N_VDD_XI9.XI172.MM4_s N_VDD_XI9.XI103.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=5.4375e-13 AS=7.65e-13 PD=7.25e-07 PS=2.52e-06
mXI9.XI171.MM4 N_XI9.XI171.NET25_XI9.XI171.MM4_d N_XI9.NET72_XI9.XI171.MM4_g
+ N_VDD_XI9.XI171.MM4_s N_VDD_XI9.XI102.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=5.4375e-13 AS=7.65e-13 PD=7.25e-07 PS=2.52e-06
mXI9.XI170.MM4 N_XI9.XI170.NET25_XI9.XI170.MM4_d N_XI9.NET60_XI9.XI170.MM4_g
+ N_VDD_XI9.XI170.MM4_s N_VDD_XI9.XI88.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=5.4375e-13 AS=7.65e-13 PD=7.25e-07 PS=2.52e-06
mXI9.XI96.MM4 N_XI9.XI96.NET25_XI9.XI96.MM4_d N_XI9.NET183_XI9.XI96.MM4_g
+ N_VDD_XI9.XI96.MM4_s N_VDD_XI9.XI82.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=5.4375e-13 AS=7.65e-13 PD=7.25e-07 PS=2.52e-06
mXI9.XI93.MM4 N_XI9.XI93.NET25_XI9.XI93.MM4_d N_XI9.NET178_XI9.XI93.MM4_g
+ N_VDD_XI9.XI93.MM4_s N_VDD_XI9.XI97.XI4.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=5.4375e-13 AS=7.65e-13 PD=7.25e-07 PS=2.52e-06
mXI9.XI182.XI9.MM1 N_XI9.XI182.NET43_XI9.XI182.XI9.MM1_d
+ N_XI9.P16_XI9.XI182.XI9.MM1_g N_VDD_XI9.XI182.XI9.MM1_s
+ N_VDD_XI9.XI153.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI9.XI181.XI9.MM1 N_XI9.XI181.NET43_XI9.XI181.XI9.MM1_d
+ N_XI9.P15_XI9.XI181.XI9.MM1_g N_VDD_XI9.XI181.XI9.MM1_s
+ N_VDD_XI9.XI154.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI9.XI180.XI9.MM1 N_XI9.XI180.NET43_XI9.XI180.XI9.MM1_d
+ N_XI9.P14_XI9.XI180.XI9.MM1_g N_VDD_XI9.XI180.XI9.MM1_s
+ N_VDD_XI9.XI157.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI9.XI179.XI4.MM1 N_XI9.XI179.NET39_XI9.XI179.XI4.MM1_d
+ N_XI9.P13_XI9.XI179.XI4.MM1_g N_VDD_XI9.XI179.XI4.MM1_s
+ N_VDD_XI9.XI156.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI9.XI178.XI9.MM1 N_XI9.XI178.NET43_XI9.XI178.XI9.MM1_d
+ N_XI9.P12_XI9.XI178.XI9.MM1_g N_VDD_XI9.XI178.XI9.MM1_s
+ N_VDD_XI9.XI155.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI9.XI177.XI9.MM1 N_XI9.XI177.NET43_XI9.XI177.XI9.MM1_d
+ N_XI9.P11_XI9.XI177.XI9.MM1_g N_VDD_XI9.XI177.XI9.MM1_s
+ N_VDD_XI9.XI133.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI9.XI176.XI9.MM1 N_XI9.XI176.NET43_XI9.XI176.XI9.MM1_d
+ N_XI9.P10_XI9.XI176.XI9.MM1_g N_VDD_XI9.XI176.XI9.MM1_s
+ N_VDD_XI9.XI132.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI9.XI175.XI9.MM1 N_XI9.XI175.NET43_XI9.XI175.XI9.MM1_d
+ N_XI9.P9_XI9.XI175.XI9.MM1_g N_VDD_XI9.XI175.XI9.MM1_s
+ N_VDD_XI9.XI131.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI9.XI174.XI9.MM1 N_XI9.XI174.NET43_XI9.XI174.XI9.MM1_d
+ N_XI9.P8_XI9.XI174.XI9.MM1_g N_VDD_XI9.XI174.XI9.MM1_s
+ N_VDD_XI9.XI111.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI9.XI173.XI9.MM1 N_XI9.XI173.NET43_XI9.XI173.XI9.MM1_d
+ N_XI9.P7_XI9.XI173.XI9.MM1_g N_VDD_XI9.XI173.XI9.MM1_s
+ N_VDD_XI9.XI110.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI9.XI172.XI9.MM1 N_XI9.XI172.NET43_XI9.XI172.XI9.MM1_d
+ N_XI9.P6_XI9.XI172.XI9.MM1_g N_VDD_XI9.XI172.XI9.MM1_s
+ N_VDD_XI9.XI103.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI9.XI171.XI9.MM1 N_XI9.XI171.NET43_XI9.XI171.XI9.MM1_d
+ N_XI9.P5_XI9.XI171.XI9.MM1_g N_VDD_XI9.XI171.XI9.MM1_s
+ N_VDD_XI9.XI102.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI9.XI170.XI9.MM1 N_XI9.XI170.NET43_XI9.XI170.XI9.MM1_d
+ N_XI9.P4_XI9.XI170.XI9.MM1_g N_VDD_XI9.XI170.XI9.MM1_s
+ N_VDD_XI9.XI88.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI9.XI96.XI9.MM1 N_XI9.XI96.NET43_XI9.XI96.XI9.MM1_d
+ N_XI9.P3_XI9.XI96.XI9.MM1_g N_VDD_XI9.XI96.XI9.MM1_s N_VDD_XI9.XI82.XI1.MM1_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI9.XI93.XI9.MM1 N_XI9.XI93.NET43_XI9.XI93.XI9.MM1_d
+ N_XI9.P2_XI9.XI93.XI9.MM1_g N_VDD_XI9.XI93.XI9.MM1_s N_VDD_XI9.XI97.XI4.MM1_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI16.XI30.XI1.MM1 N_XI16.XI30.NET6_XI16.XI30.XI1.MM1_d
+ N_NET198_XI16.XI30.XI1.MM1_g N_VDD_XI16.XI30.XI1.MM1_s
+ N_VDD_XI16.XI30.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=4.125e-13 AS=7.35e-13
+ PD=5.5e-07 PS=2.48e-06
mXI16.XI29.XI1.MM1 N_XI16.XI29.NET6_XI16.XI29.XI1.MM1_d
+ N_NET198_XI16.XI29.XI1.MM1_g N_VDD_XI16.XI29.XI1.MM1_s
+ N_VDD_XI16.XI29.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=4.125e-13 AS=7.35e-13
+ PD=5.5e-07 PS=2.48e-06
mXI16.XI28.XI1.MM1 N_XI16.XI28.NET6_XI16.XI28.XI1.MM1_d
+ N_NET198_XI16.XI28.XI1.MM1_g N_VDD_XI16.XI28.XI1.MM1_s
+ N_VDD_XI16.XI28.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=4.125e-13 AS=7.35e-13
+ PD=5.5e-07 PS=2.48e-06
mXI16.XI27.XI1.MM1 N_XI16.XI27.NET6_XI16.XI27.XI1.MM1_d
+ N_NET198_XI16.XI27.XI1.MM1_g N_VDD_XI16.XI27.XI1.MM1_s
+ N_VDD_XI16.XI27.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=4.125e-13 AS=7.35e-13
+ PD=5.5e-07 PS=2.48e-06
mXI16.XI26.XI1.MM1 N_XI16.XI26.NET6_XI16.XI26.XI1.MM1_d
+ N_NET198_XI16.XI26.XI1.MM1_g N_VDD_XI16.XI26.XI1.MM1_s
+ N_VDD_XI16.XI26.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=4.125e-13 AS=7.35e-13
+ PD=5.5e-07 PS=2.48e-06
mXI16.XI25.XI1.MM1 N_XI16.XI25.NET6_XI16.XI25.XI1.MM1_d
+ N_NET198_XI16.XI25.XI1.MM1_g N_VDD_XI16.XI25.XI1.MM1_s
+ N_VDD_XI16.XI25.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=4.125e-13 AS=7.35e-13
+ PD=5.5e-07 PS=2.48e-06
mXI16.XI24.XI1.MM1 N_XI16.XI24.NET6_XI16.XI24.XI1.MM1_d
+ N_NET198_XI16.XI24.XI1.MM1_g N_VDD_XI16.XI24.XI1.MM1_s
+ N_VDD_XI16.XI24.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=4.125e-13 AS=7.35e-13
+ PD=5.5e-07 PS=2.48e-06
mXI16.XI23.XI1.MM1 N_XI16.XI23.NET6_XI16.XI23.XI1.MM1_d
+ N_NET198_XI16.XI23.XI1.MM1_g N_VDD_XI16.XI23.XI1.MM1_s
+ N_VDD_XI16.XI23.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=4.125e-13 AS=7.35e-13
+ PD=5.5e-07 PS=2.48e-06
mXI16.XI22.XI1.MM1 N_XI16.XI22.NET6_XI16.XI22.XI1.MM1_d
+ N_NET198_XI16.XI22.XI1.MM1_g N_VDD_XI16.XI22.XI1.MM1_s
+ N_VDD_XI16.XI22.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=4.125e-13 AS=7.35e-13
+ PD=5.5e-07 PS=2.48e-06
mXI16.XI21.XI1.MM1 N_XI16.XI21.NET6_XI16.XI21.XI1.MM1_d
+ N_NET198_XI16.XI21.XI1.MM1_g N_VDD_XI16.XI21.XI1.MM1_s
+ N_VDD_XI16.XI21.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=4.125e-13 AS=7.35e-13
+ PD=5.5e-07 PS=2.48e-06
mXI16.XI20.XI1.MM1 N_XI16.XI20.NET6_XI16.XI20.XI1.MM1_d
+ N_NET198_XI16.XI20.XI1.MM1_g N_VDD_XI16.XI20.XI1.MM1_s
+ N_VDD_XI16.XI20.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=4.125e-13 AS=7.35e-13
+ PD=5.5e-07 PS=2.48e-06
mXI16.XI19.XI1.MM1 N_XI16.XI19.NET6_XI16.XI19.XI1.MM1_d
+ N_NET198_XI16.XI19.XI1.MM1_g N_VDD_XI16.XI19.XI1.MM1_s
+ N_VDD_XI16.XI19.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=4.125e-13 AS=7.35e-13
+ PD=5.5e-07 PS=2.48e-06
mXI16.XI18.XI1.MM1 N_XI16.XI18.NET6_XI16.XI18.XI1.MM1_d
+ N_NET198_XI16.XI18.XI1.MM1_g N_VDD_XI16.XI18.XI1.MM1_s
+ N_VDD_XI16.XI18.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=4.125e-13 AS=7.35e-13
+ PD=5.5e-07 PS=2.48e-06
mXI16.XI17.XI1.MM1 N_XI16.XI17.NET6_XI16.XI17.XI1.MM1_d
+ N_NET198_XI16.XI17.XI1.MM1_g N_VDD_XI16.XI17.XI1.MM1_s
+ N_VDD_XI16.XI17.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=4.125e-13 AS=7.35e-13
+ PD=5.5e-07 PS=2.48e-06
mXI16.XI16.XI1.MM1 N_XI16.XI16.NET6_XI16.XI16.XI1.MM1_d
+ N_NET198_XI16.XI16.XI1.MM1_g N_VDD_XI16.XI16.XI1.MM1_s
+ N_VDD_XI16.XI16.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=4.125e-13 AS=7.35e-13
+ PD=5.5e-07 PS=2.48e-06
mXI16.XI0.XI1.MM3 N_XI16.XI0.NET6_XI16.XI0.XI1.MM3_d N_NET198_XI16.XI0.XI1.MM3_g
+ N_VDD_XI16.XI0.XI1.MM3_s N_VDD_XI16.XI0.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=4.125e-13 AS=7.35e-13 PD=5.5e-07 PS=2.48e-06
mXI16.XI30.XI1.MM3 N_XI16.XI30.NET6_XI16.XI30.XI1.MM3_d
+ N_NET177_XI16.XI30.XI1.MM3_g N_VDD_XI16.XI30.XI1.MM3_s
+ N_VDD_XI16.XI30.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=4.125e-13 AS=7.65e-13
+ PD=5.5e-07 PS=2.52e-06
mXI16.XI29.XI1.MM3 N_XI16.XI29.NET6_XI16.XI29.XI1.MM3_d
+ N_NET178_XI16.XI29.XI1.MM3_g N_VDD_XI16.XI29.XI1.MM3_s
+ N_VDD_XI16.XI29.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=4.125e-13 AS=7.65e-13
+ PD=5.5e-07 PS=2.52e-06
mXI16.XI28.XI1.MM3 N_XI16.XI28.NET6_XI16.XI28.XI1.MM3_d
+ N_NET179_XI16.XI28.XI1.MM3_g N_VDD_XI16.XI28.XI1.MM3_s
+ N_VDD_XI16.XI28.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=4.125e-13 AS=7.65e-13
+ PD=5.5e-07 PS=2.52e-06
mXI16.XI27.XI1.MM3 N_XI16.XI27.NET6_XI16.XI27.XI1.MM3_d
+ N_NET180_XI16.XI27.XI1.MM3_g N_VDD_XI16.XI27.XI1.MM3_s
+ N_VDD_XI16.XI27.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=4.125e-13 AS=7.65e-13
+ PD=5.5e-07 PS=2.52e-06
mXI16.XI26.XI1.MM3 N_XI16.XI26.NET6_XI16.XI26.XI1.MM3_d
+ N_NET181_XI16.XI26.XI1.MM3_g N_VDD_XI16.XI26.XI1.MM3_s
+ N_VDD_XI16.XI26.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=4.125e-13 AS=7.65e-13
+ PD=5.5e-07 PS=2.52e-06
mXI16.XI25.XI1.MM3 N_XI16.XI25.NET6_XI16.XI25.XI1.MM3_d
+ N_NET182_XI16.XI25.XI1.MM3_g N_VDD_XI16.XI25.XI1.MM3_s
+ N_VDD_XI16.XI25.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=4.125e-13 AS=7.65e-13
+ PD=5.5e-07 PS=2.52e-06
mXI16.XI24.XI1.MM3 N_XI16.XI24.NET6_XI16.XI24.XI1.MM3_d
+ N_NET183_XI16.XI24.XI1.MM3_g N_VDD_XI16.XI24.XI1.MM3_s
+ N_VDD_XI16.XI24.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=4.125e-13 AS=7.65e-13
+ PD=5.5e-07 PS=2.52e-06
mXI16.XI23.XI1.MM3 N_XI16.XI23.NET6_XI16.XI23.XI1.MM3_d
+ N_NET184_XI16.XI23.XI1.MM3_g N_VDD_XI16.XI23.XI1.MM3_s
+ N_VDD_XI16.XI23.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=4.125e-13 AS=7.65e-13
+ PD=5.5e-07 PS=2.52e-06
mXI16.XI22.XI1.MM3 N_XI16.XI22.NET6_XI16.XI22.XI1.MM3_d
+ N_NET185_XI16.XI22.XI1.MM3_g N_VDD_XI16.XI22.XI1.MM3_s
+ N_VDD_XI16.XI22.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=4.125e-13 AS=7.65e-13
+ PD=5.5e-07 PS=2.52e-06
mXI16.XI21.XI1.MM3 N_XI16.XI21.NET6_XI16.XI21.XI1.MM3_d
+ N_NET186_XI16.XI21.XI1.MM3_g N_VDD_XI16.XI21.XI1.MM3_s
+ N_VDD_XI16.XI21.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=4.125e-13 AS=7.65e-13
+ PD=5.5e-07 PS=2.52e-06
mXI16.XI20.XI1.MM3 N_XI16.XI20.NET6_XI16.XI20.XI1.MM3_d
+ N_NET187_XI16.XI20.XI1.MM3_g N_VDD_XI16.XI20.XI1.MM3_s
+ N_VDD_XI16.XI20.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=4.125e-13 AS=7.65e-13
+ PD=5.5e-07 PS=2.52e-06
mXI16.XI19.XI1.MM3 N_XI16.XI19.NET6_XI16.XI19.XI1.MM3_d
+ N_NET188_XI16.XI19.XI1.MM3_g N_VDD_XI16.XI19.XI1.MM3_s
+ N_VDD_XI16.XI19.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=4.125e-13 AS=7.65e-13
+ PD=5.5e-07 PS=2.52e-06
mXI16.XI18.XI1.MM3 N_XI16.XI18.NET6_XI16.XI18.XI1.MM3_d
+ N_NET189_XI16.XI18.XI1.MM3_g N_VDD_XI16.XI18.XI1.MM3_s
+ N_VDD_XI16.XI18.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=4.125e-13 AS=7.65e-13
+ PD=5.5e-07 PS=2.52e-06
mXI16.XI17.XI1.MM3 N_XI16.XI17.NET6_XI16.XI17.XI1.MM3_d
+ N_NET190_XI16.XI17.XI1.MM3_g N_VDD_XI16.XI17.XI1.MM3_s
+ N_VDD_XI16.XI17.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=4.125e-13 AS=7.65e-13
+ PD=5.5e-07 PS=2.52e-06
mXI16.XI16.XI1.MM3 N_XI16.XI16.NET6_XI16.XI16.XI1.MM3_d
+ N_NET191_XI16.XI16.XI1.MM3_g N_VDD_XI16.XI16.XI1.MM3_s
+ N_VDD_XI16.XI16.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=4.125e-13 AS=7.65e-13
+ PD=5.5e-07 PS=2.52e-06
mXI16.XI0.XI1.MM1 N_XI16.XI0.NET6_XI16.XI0.XI1.MM1_d N_NET192_XI16.XI0.XI1.MM1_g
+ N_VDD_XI16.XI0.XI1.MM1_s N_VDD_XI16.XI0.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=4.125e-13 AS=7.65e-13 PD=5.5e-07 PS=2.52e-06
mXI16.XI30.XI0.MM1 N_NET452_XI16.XI30.XI0.MM1_d
+ N_XI16.XI30.NET6_XI16.XI30.XI0.MM1_g N_VDD_XI16.XI30.XI0.MM1_s
+ N_VDD_XI16.XI30.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI16.XI29.XI0.MM1 N_NET453_XI16.XI29.XI0.MM1_d
+ N_XI16.XI29.NET6_XI16.XI29.XI0.MM1_g N_VDD_XI16.XI29.XI0.MM1_s
+ N_VDD_XI16.XI29.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI16.XI28.XI0.MM1 N_NET454_XI16.XI28.XI0.MM1_d
+ N_XI16.XI28.NET6_XI16.XI28.XI0.MM1_g N_VDD_XI16.XI28.XI0.MM1_s
+ N_VDD_XI16.XI28.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI16.XI27.XI0.MM1 N_NET455_XI16.XI27.XI0.MM1_d
+ N_XI16.XI27.NET6_XI16.XI27.XI0.MM1_g N_VDD_XI16.XI27.XI0.MM1_s
+ N_VDD_XI16.XI27.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI16.XI26.XI0.MM1 N_NET456_XI16.XI26.XI0.MM1_d
+ N_XI16.XI26.NET6_XI16.XI26.XI0.MM1_g N_VDD_XI16.XI26.XI0.MM1_s
+ N_VDD_XI16.XI26.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI16.XI25.XI0.MM1 N_NET457_XI16.XI25.XI0.MM1_d
+ N_XI16.XI25.NET6_XI16.XI25.XI0.MM1_g N_VDD_XI16.XI25.XI0.MM1_s
+ N_VDD_XI16.XI25.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI16.XI24.XI0.MM1 N_NET458_XI16.XI24.XI0.MM1_d
+ N_XI16.XI24.NET6_XI16.XI24.XI0.MM1_g N_VDD_XI16.XI24.XI0.MM1_s
+ N_VDD_XI16.XI24.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI16.XI23.XI0.MM1 N_NET459_XI16.XI23.XI0.MM1_d
+ N_XI16.XI23.NET6_XI16.XI23.XI0.MM1_g N_VDD_XI16.XI23.XI0.MM1_s
+ N_VDD_XI16.XI23.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI16.XI22.XI0.MM1 N_NET460_XI16.XI22.XI0.MM1_d
+ N_XI16.XI22.NET6_XI16.XI22.XI0.MM1_g N_VDD_XI16.XI22.XI0.MM1_s
+ N_VDD_XI16.XI22.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI16.XI21.XI0.MM1 N_NET461_XI16.XI21.XI0.MM1_d
+ N_XI16.XI21.NET6_XI16.XI21.XI0.MM1_g N_VDD_XI16.XI21.XI0.MM1_s
+ N_VDD_XI16.XI21.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI16.XI20.XI0.MM1 N_NET462_XI16.XI20.XI0.MM1_d
+ N_XI16.XI20.NET6_XI16.XI20.XI0.MM1_g N_VDD_XI16.XI20.XI0.MM1_s
+ N_VDD_XI16.XI20.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI16.XI19.XI0.MM1 N_NET463_XI16.XI19.XI0.MM1_d
+ N_XI16.XI19.NET6_XI16.XI19.XI0.MM1_g N_VDD_XI16.XI19.XI0.MM1_s
+ N_VDD_XI16.XI19.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI16.XI18.XI0.MM1 N_NET464_XI16.XI18.XI0.MM1_d
+ N_XI16.XI18.NET6_XI16.XI18.XI0.MM1_g N_VDD_XI16.XI18.XI0.MM1_s
+ N_VDD_XI16.XI18.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI16.XI17.XI0.MM1 N_NET465_XI16.XI17.XI0.MM1_d
+ N_XI16.XI17.NET6_XI16.XI17.XI0.MM1_g N_VDD_XI16.XI17.XI0.MM1_s
+ N_VDD_XI16.XI17.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI16.XI16.XI0.MM1 N_NET466_XI16.XI16.XI0.MM1_d
+ N_XI16.XI16.NET6_XI16.XI16.XI0.MM1_g N_VDD_XI16.XI16.XI0.MM1_s
+ N_VDD_XI16.XI16.XI1.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI16.XI0.XI0.MM1 N_NET467_XI16.XI0.XI0.MM1_d N_XI16.XI0.NET6_XI16.XI0.XI0.MM1_g
+ N_VDD_XI16.XI0.XI0.MM1_s N_VDD_XI16.XI0.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI11.XI30.XI0.MM1 N_XI11.XI30.NET0180_XI11.XI30.XI0.MM1_d
+ N_NET222_XI11.XI30.XI0.MM1_g N_VDD_XI11.XI30.XI0.MM1_s
+ N_VDD_XI11.XI30.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI11.XI29.XI0.MM1 N_XI11.XI29.NET0180_XI11.XI29.XI0.MM1_d
+ N_NET222_XI11.XI29.XI0.MM1_g N_VDD_XI11.XI29.XI0.MM1_s
+ N_VDD_XI11.XI29.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI11.XI31.XI0.MM1 N_XI11.XI31.NET0180_XI11.XI31.XI0.MM1_d
+ N_NET222_XI11.XI31.XI0.MM1_g N_VDD_XI11.XI31.XI0.MM1_s
+ N_VDD_XI11.XI31.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI11.XI28.XI0.MM1 N_XI11.XI28.NET0180_XI11.XI28.XI0.MM1_d
+ N_NET222_XI11.XI28.XI0.MM1_g N_VDD_XI11.XI28.XI0.MM1_s
+ N_VDD_XI11.XI28.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI11.XI25.XI0.MM1 N_XI11.XI25.NET0180_XI11.XI25.XI0.MM1_d
+ N_NET222_XI11.XI25.XI0.MM1_g N_VDD_XI11.XI25.XI0.MM1_s
+ N_VDD_XI11.XI25.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI11.XI26.XI0.MM1 N_XI11.XI26.NET0180_XI11.XI26.XI0.MM1_d
+ N_NET222_XI11.XI26.XI0.MM1_g N_VDD_XI11.XI26.XI0.MM1_s
+ N_VDD_XI11.XI26.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI11.XI24.XI0.MM1 N_XI11.XI24.NET0180_XI11.XI24.XI0.MM1_d
+ N_NET222_XI11.XI24.XI0.MM1_g N_VDD_XI11.XI24.XI0.MM1_s
+ N_VDD_XI11.XI24.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI11.XI27.XI0.MM1 N_XI11.XI27.NET0180_XI11.XI27.XI0.MM1_d
+ N_NET222_XI11.XI27.XI0.MM1_g N_VDD_XI11.XI27.XI0.MM1_s
+ N_VDD_XI11.XI27.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI11.XI22.XI0.MM1 N_XI11.XI22.NET0180_XI11.XI22.XI0.MM1_d
+ N_NET222_XI11.XI22.XI0.MM1_g N_VDD_XI11.XI22.XI0.MM1_s
+ N_VDD_XI11.XI22.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI11.XI21.XI0.MM1 N_XI11.XI21.NET0180_XI11.XI21.XI0.MM1_d
+ N_NET222_XI11.XI21.XI0.MM1_g N_VDD_XI11.XI21.XI0.MM1_s
+ N_VDD_XI11.XI21.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI11.XI23.XI0.MM1 N_XI11.XI23.NET0180_XI11.XI23.XI0.MM1_d
+ N_NET222_XI11.XI23.XI0.MM1_g N_VDD_XI11.XI23.XI0.MM1_s
+ N_VDD_XI11.XI23.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI11.XI19.XI0.MM1 N_XI11.XI19.NET0180_XI11.XI19.XI0.MM1_d
+ N_NET222_XI11.XI19.XI0.MM1_g N_VDD_XI11.XI19.XI0.MM1_s
+ N_VDD_XI11.XI19.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI11.XI20.XI0.MM1 N_XI11.XI20.NET0180_XI11.XI20.XI0.MM1_d
+ N_NET222_XI11.XI20.XI0.MM1_g N_VDD_XI11.XI20.XI0.MM1_s
+ N_VDD_XI11.XI20.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI11.XI18.XI0.MM1 N_XI11.XI18.NET0180_XI11.XI18.XI0.MM1_d
+ N_NET222_XI11.XI18.XI0.MM1_g N_VDD_XI11.XI18.XI0.MM1_s
+ N_VDD_XI11.XI18.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI11.XI17.XI0.MM1 N_XI11.XI17.NET0180_XI11.XI17.XI0.MM1_d
+ N_NET222_XI11.XI17.XI0.MM1_g N_VDD_XI11.XI17.XI0.MM1_s
+ N_VDD_XI11.XI17.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI11.XI0.XI0.MM1 N_XI11.XI0.NET0180_XI11.XI0.XI0.MM1_d
+ N_NET222_XI11.XI0.XI0.MM1_g N_VDD_XI11.XI0.XI0.MM1_s N_VDD_XI11.XI0.XI0.MM1_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI11.XI30.XI1.MM1 N_XI11.XI30.NET35_XI11.XI30.XI1.MM1_d
+ N_XI11.XI30.NET0180_XI11.XI30.XI1.MM1_g N_VDD_XI11.XI30.XI1.MM1_s
+ N_VDD_XI11.XI30.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI11.XI29.XI1.MM1 N_XI11.XI29.NET35_XI11.XI29.XI1.MM1_d
+ N_XI11.XI29.NET0180_XI11.XI29.XI1.MM1_g N_VDD_XI11.XI29.XI1.MM1_s
+ N_VDD_XI11.XI29.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI11.XI31.XI1.MM1 N_XI11.XI31.NET35_XI11.XI31.XI1.MM1_d
+ N_XI11.XI31.NET0180_XI11.XI31.XI1.MM1_g N_VDD_XI11.XI31.XI1.MM1_s
+ N_VDD_XI11.XI31.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI11.XI28.XI1.MM1 N_XI11.XI28.NET35_XI11.XI28.XI1.MM1_d
+ N_XI11.XI28.NET0180_XI11.XI28.XI1.MM1_g N_VDD_XI11.XI28.XI1.MM1_s
+ N_VDD_XI11.XI28.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI11.XI25.XI1.MM1 N_XI11.XI25.NET35_XI11.XI25.XI1.MM1_d
+ N_XI11.XI25.NET0180_XI11.XI25.XI1.MM1_g N_VDD_XI11.XI25.XI1.MM1_s
+ N_VDD_XI11.XI25.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI11.XI26.XI1.MM1 N_XI11.XI26.NET35_XI11.XI26.XI1.MM1_d
+ N_XI11.XI26.NET0180_XI11.XI26.XI1.MM1_g N_VDD_XI11.XI26.XI1.MM1_s
+ N_VDD_XI11.XI26.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI11.XI24.XI1.MM1 N_XI11.XI24.NET35_XI11.XI24.XI1.MM1_d
+ N_XI11.XI24.NET0180_XI11.XI24.XI1.MM1_g N_VDD_XI11.XI24.XI1.MM1_s
+ N_VDD_XI11.XI24.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI11.XI27.XI1.MM1 N_XI11.XI27.NET35_XI11.XI27.XI1.MM1_d
+ N_XI11.XI27.NET0180_XI11.XI27.XI1.MM1_g N_VDD_XI11.XI27.XI1.MM1_s
+ N_VDD_XI11.XI27.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI11.XI22.XI1.MM1 N_XI11.XI22.NET35_XI11.XI22.XI1.MM1_d
+ N_XI11.XI22.NET0180_XI11.XI22.XI1.MM1_g N_VDD_XI11.XI22.XI1.MM1_s
+ N_VDD_XI11.XI22.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI11.XI21.XI1.MM1 N_XI11.XI21.NET35_XI11.XI21.XI1.MM1_d
+ N_XI11.XI21.NET0180_XI11.XI21.XI1.MM1_g N_VDD_XI11.XI21.XI1.MM1_s
+ N_VDD_XI11.XI21.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI11.XI23.XI1.MM1 N_XI11.XI23.NET35_XI11.XI23.XI1.MM1_d
+ N_XI11.XI23.NET0180_XI11.XI23.XI1.MM1_g N_VDD_XI11.XI23.XI1.MM1_s
+ N_VDD_XI11.XI23.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI11.XI19.XI1.MM1 N_XI11.XI19.NET35_XI11.XI19.XI1.MM1_d
+ N_XI11.XI19.NET0180_XI11.XI19.XI1.MM1_g N_VDD_XI11.XI19.XI1.MM1_s
+ N_VDD_XI11.XI19.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI11.XI20.XI1.MM1 N_XI11.XI20.NET35_XI11.XI20.XI1.MM1_d
+ N_XI11.XI20.NET0180_XI11.XI20.XI1.MM1_g N_VDD_XI11.XI20.XI1.MM1_s
+ N_VDD_XI11.XI20.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI11.XI18.XI1.MM1 N_XI11.XI18.NET35_XI11.XI18.XI1.MM1_d
+ N_XI11.XI18.NET0180_XI11.XI18.XI1.MM1_g N_VDD_XI11.XI18.XI1.MM1_s
+ N_VDD_XI11.XI18.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI11.XI17.XI1.MM1 N_XI11.XI17.NET35_XI11.XI17.XI1.MM1_d
+ N_XI11.XI17.NET0180_XI11.XI17.XI1.MM1_g N_VDD_XI11.XI17.XI1.MM1_s
+ N_VDD_XI11.XI17.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI11.XI0.XI1.MM1 N_XI11.XI0.NET35_XI11.XI0.XI1.MM1_d
+ N_XI11.XI0.NET0180_XI11.XI0.XI1.MM1_g N_VDD_XI11.XI0.XI1.MM1_s
+ N_VDD_XI11.XI0.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI11.XI30.MM25 N_XI11.XI30.CLKB_XI11.XI30.MM25_d
+ N_XI11.XI30.NET35_XI11.XI30.MM25_g N_VDD_XI11.XI30.MM25_s
+ N_VDD_XI11.XI30.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI11.XI29.MM25 N_XI11.XI29.CLKB_XI11.XI29.MM25_d
+ N_XI11.XI29.NET35_XI11.XI29.MM25_g N_VDD_XI11.XI29.MM25_s
+ N_VDD_XI11.XI29.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI11.XI31.MM25 N_XI11.XI31.CLKB_XI11.XI31.MM25_d
+ N_XI11.XI31.NET35_XI11.XI31.MM25_g N_VDD_XI11.XI31.MM25_s
+ N_VDD_XI11.XI31.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI11.XI28.MM25 N_XI11.XI28.CLKB_XI11.XI28.MM25_d
+ N_XI11.XI28.NET35_XI11.XI28.MM25_g N_VDD_XI11.XI28.MM25_s
+ N_VDD_XI11.XI28.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI11.XI25.MM25 N_XI11.XI25.CLKB_XI11.XI25.MM25_d
+ N_XI11.XI25.NET35_XI11.XI25.MM25_g N_VDD_XI11.XI25.MM25_s
+ N_VDD_XI11.XI25.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI11.XI26.MM25 N_XI11.XI26.CLKB_XI11.XI26.MM25_d
+ N_XI11.XI26.NET35_XI11.XI26.MM25_g N_VDD_XI11.XI26.MM25_s
+ N_VDD_XI11.XI26.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI11.XI24.MM25 N_XI11.XI24.CLKB_XI11.XI24.MM25_d
+ N_XI11.XI24.NET35_XI11.XI24.MM25_g N_VDD_XI11.XI24.MM25_s
+ N_VDD_XI11.XI24.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI11.XI27.MM25 N_XI11.XI27.CLKB_XI11.XI27.MM25_d
+ N_XI11.XI27.NET35_XI11.XI27.MM25_g N_VDD_XI11.XI27.MM25_s
+ N_VDD_XI11.XI27.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI11.XI22.MM25 N_XI11.XI22.CLKB_XI11.XI22.MM25_d
+ N_XI11.XI22.NET35_XI11.XI22.MM25_g N_VDD_XI11.XI22.MM25_s
+ N_VDD_XI11.XI22.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI11.XI21.MM25 N_XI11.XI21.CLKB_XI11.XI21.MM25_d
+ N_XI11.XI21.NET35_XI11.XI21.MM25_g N_VDD_XI11.XI21.MM25_s
+ N_VDD_XI11.XI21.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI11.XI23.MM25 N_XI11.XI23.CLKB_XI11.XI23.MM25_d
+ N_XI11.XI23.NET35_XI11.XI23.MM25_g N_VDD_XI11.XI23.MM25_s
+ N_VDD_XI11.XI23.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI11.XI19.MM25 N_XI11.XI19.CLKB_XI11.XI19.MM25_d
+ N_XI11.XI19.NET35_XI11.XI19.MM25_g N_VDD_XI11.XI19.MM25_s
+ N_VDD_XI11.XI19.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI11.XI20.MM25 N_XI11.XI20.CLKB_XI11.XI20.MM25_d
+ N_XI11.XI20.NET35_XI11.XI20.MM25_g N_VDD_XI11.XI20.MM25_s
+ N_VDD_XI11.XI20.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI11.XI18.MM25 N_XI11.XI18.CLKB_XI11.XI18.MM25_d
+ N_XI11.XI18.NET35_XI11.XI18.MM25_g N_VDD_XI11.XI18.MM25_s
+ N_VDD_XI11.XI18.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI11.XI17.MM25 N_XI11.XI17.CLKB_XI11.XI17.MM25_d
+ N_XI11.XI17.NET35_XI11.XI17.MM25_g N_VDD_XI11.XI17.MM25_s
+ N_VDD_XI11.XI17.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI11.XI0.MM25 N_XI11.XI0.CLKB_XI11.XI0.MM25_d N_XI11.XI0.NET35_XI11.XI0.MM25_g
+ N_VDD_XI11.XI0.MM25_s N_VDD_XI11.XI0.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI11.XI30.MM20 N_XI11.XI30.NET27_XI11.XI30.MM20_d N_NET452_XI11.XI30.MM20_g
+ N_VDD_XI11.XI30.MM20_s N_VDD_XI11.XI30.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI11.XI29.MM20 N_XI11.XI29.NET27_XI11.XI29.MM20_d N_NET453_XI11.XI29.MM20_g
+ N_VDD_XI11.XI29.MM20_s N_VDD_XI11.XI29.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI11.XI31.MM20 N_XI11.XI31.NET27_XI11.XI31.MM20_d N_NET454_XI11.XI31.MM20_g
+ N_VDD_XI11.XI31.MM20_s N_VDD_XI11.XI31.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI11.XI28.MM20 N_XI11.XI28.NET27_XI11.XI28.MM20_d N_NET455_XI11.XI28.MM20_g
+ N_VDD_XI11.XI28.MM20_s N_VDD_XI11.XI28.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI11.XI25.MM20 N_XI11.XI25.NET27_XI11.XI25.MM20_d N_NET456_XI11.XI25.MM20_g
+ N_VDD_XI11.XI25.MM20_s N_VDD_XI11.XI25.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI11.XI26.MM20 N_XI11.XI26.NET27_XI11.XI26.MM20_d N_NET457_XI11.XI26.MM20_g
+ N_VDD_XI11.XI26.MM20_s N_VDD_XI11.XI26.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI11.XI24.MM20 N_XI11.XI24.NET27_XI11.XI24.MM20_d N_NET458_XI11.XI24.MM20_g
+ N_VDD_XI11.XI24.MM20_s N_VDD_XI11.XI24.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI11.XI27.MM20 N_XI11.XI27.NET27_XI11.XI27.MM20_d N_NET459_XI11.XI27.MM20_g
+ N_VDD_XI11.XI27.MM20_s N_VDD_XI11.XI27.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI11.XI22.MM20 N_XI11.XI22.NET27_XI11.XI22.MM20_d N_NET460_XI11.XI22.MM20_g
+ N_VDD_XI11.XI22.MM20_s N_VDD_XI11.XI22.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI11.XI21.MM20 N_XI11.XI21.NET27_XI11.XI21.MM20_d N_NET461_XI11.XI21.MM20_g
+ N_VDD_XI11.XI21.MM20_s N_VDD_XI11.XI21.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI11.XI23.MM20 N_XI11.XI23.NET27_XI11.XI23.MM20_d N_NET462_XI11.XI23.MM20_g
+ N_VDD_XI11.XI23.MM20_s N_VDD_XI11.XI23.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI11.XI19.MM20 N_XI11.XI19.NET27_XI11.XI19.MM20_d N_NET463_XI11.XI19.MM20_g
+ N_VDD_XI11.XI19.MM20_s N_VDD_XI11.XI19.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI11.XI20.MM20 N_XI11.XI20.NET27_XI11.XI20.MM20_d N_NET464_XI11.XI20.MM20_g
+ N_VDD_XI11.XI20.MM20_s N_VDD_XI11.XI20.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI11.XI18.MM20 N_XI11.XI18.NET27_XI11.XI18.MM20_d N_NET465_XI11.XI18.MM20_g
+ N_VDD_XI11.XI18.MM20_s N_VDD_XI11.XI18.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI11.XI17.MM20 N_XI11.XI17.NET27_XI11.XI17.MM20_d N_NET466_XI11.XI17.MM20_g
+ N_VDD_XI11.XI17.MM20_s N_VDD_XI11.XI17.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI11.XI0.MM20 N_XI11.XI0.NET27_XI11.XI0.MM20_d N_NET467_XI11.XI0.MM20_g
+ N_VDD_XI11.XI0.MM20_s N_VDD_XI11.XI0.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI11.XI30.MM17 N_XI11.XI30.NET31_XI11.XI30.MM17_d
+ N_XI11.XI30.NET27_XI11.XI30.MM17_g N_VDD_XI11.XI30.MM17_s
+ N_VDD_XI11.XI30.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI11.XI29.MM17 N_XI11.XI29.NET31_XI11.XI29.MM17_d
+ N_XI11.XI29.NET27_XI11.XI29.MM17_g N_VDD_XI11.XI29.MM17_s
+ N_VDD_XI11.XI29.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI11.XI31.MM17 N_XI11.XI31.NET31_XI11.XI31.MM17_d
+ N_XI11.XI31.NET27_XI11.XI31.MM17_g N_VDD_XI11.XI31.MM17_s
+ N_VDD_XI11.XI31.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI11.XI28.MM17 N_XI11.XI28.NET31_XI11.XI28.MM17_d
+ N_XI11.XI28.NET27_XI11.XI28.MM17_g N_VDD_XI11.XI28.MM17_s
+ N_VDD_XI11.XI28.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI11.XI25.MM17 N_XI11.XI25.NET31_XI11.XI25.MM17_d
+ N_XI11.XI25.NET27_XI11.XI25.MM17_g N_VDD_XI11.XI25.MM17_s
+ N_VDD_XI11.XI25.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI11.XI26.MM17 N_XI11.XI26.NET31_XI11.XI26.MM17_d
+ N_XI11.XI26.NET27_XI11.XI26.MM17_g N_VDD_XI11.XI26.MM17_s
+ N_VDD_XI11.XI26.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI11.XI24.MM17 N_XI11.XI24.NET31_XI11.XI24.MM17_d
+ N_XI11.XI24.NET27_XI11.XI24.MM17_g N_VDD_XI11.XI24.MM17_s
+ N_VDD_XI11.XI24.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI11.XI27.MM17 N_XI11.XI27.NET31_XI11.XI27.MM17_d
+ N_XI11.XI27.NET27_XI11.XI27.MM17_g N_VDD_XI11.XI27.MM17_s
+ N_VDD_XI11.XI27.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI11.XI22.MM17 N_XI11.XI22.NET31_XI11.XI22.MM17_d
+ N_XI11.XI22.NET27_XI11.XI22.MM17_g N_VDD_XI11.XI22.MM17_s
+ N_VDD_XI11.XI22.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI11.XI21.MM17 N_XI11.XI21.NET31_XI11.XI21.MM17_d
+ N_XI11.XI21.NET27_XI11.XI21.MM17_g N_VDD_XI11.XI21.MM17_s
+ N_VDD_XI11.XI21.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI11.XI23.MM17 N_XI11.XI23.NET31_XI11.XI23.MM17_d
+ N_XI11.XI23.NET27_XI11.XI23.MM17_g N_VDD_XI11.XI23.MM17_s
+ N_VDD_XI11.XI23.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI11.XI19.MM17 N_XI11.XI19.NET31_XI11.XI19.MM17_d
+ N_XI11.XI19.NET27_XI11.XI19.MM17_g N_VDD_XI11.XI19.MM17_s
+ N_VDD_XI11.XI19.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI11.XI20.MM17 N_XI11.XI20.NET31_XI11.XI20.MM17_d
+ N_XI11.XI20.NET27_XI11.XI20.MM17_g N_VDD_XI11.XI20.MM17_s
+ N_VDD_XI11.XI20.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI11.XI18.MM17 N_XI11.XI18.NET31_XI11.XI18.MM17_d
+ N_XI11.XI18.NET27_XI11.XI18.MM17_g N_VDD_XI11.XI18.MM17_s
+ N_VDD_XI11.XI18.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI11.XI17.MM17 N_XI11.XI17.NET31_XI11.XI17.MM17_d
+ N_XI11.XI17.NET27_XI11.XI17.MM17_g N_VDD_XI11.XI17.MM17_s
+ N_VDD_XI11.XI17.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI11.XI0.MM17 N_XI11.XI0.NET31_XI11.XI0.MM17_d N_XI11.XI0.NET27_XI11.XI0.MM17_g
+ N_VDD_XI11.XI0.MM17_s N_VDD_XI11.XI0.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI11.XI30.MM27 N_XI11.XI30.NET31_XI11.XI30.MM27_d
+ N_XI11.XI30.NET35_XI11.XI30.MM27_g N_XI11.XI30.NET58_XI11.XI30.MM27_s
+ N_VDD_XI11.XI30.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=1.125e-12 AS=9.375e-13
+ PD=3e-06 PS=2.75e-06
mXI11.XI29.MM27 N_XI11.XI29.NET31_XI11.XI29.MM27_d
+ N_XI11.XI29.NET35_XI11.XI29.MM27_g N_XI11.XI29.NET58_XI11.XI29.MM27_s
+ N_VDD_XI11.XI29.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=1.125e-12 AS=9.375e-13
+ PD=3e-06 PS=2.75e-06
mXI11.XI31.MM27 N_XI11.XI31.NET31_XI11.XI31.MM27_d
+ N_XI11.XI31.NET35_XI11.XI31.MM27_g N_XI11.XI31.NET58_XI11.XI31.MM27_s
+ N_VDD_XI11.XI31.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=1.125e-12 AS=9.375e-13
+ PD=3e-06 PS=2.75e-06
mXI11.XI28.MM27 N_XI11.XI28.NET31_XI11.XI28.MM27_d
+ N_XI11.XI28.NET35_XI11.XI28.MM27_g N_XI11.XI28.NET58_XI11.XI28.MM27_s
+ N_VDD_XI11.XI28.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=1.125e-12 AS=9.375e-13
+ PD=3e-06 PS=2.75e-06
mXI11.XI25.MM27 N_XI11.XI25.NET31_XI11.XI25.MM27_d
+ N_XI11.XI25.NET35_XI11.XI25.MM27_g N_XI11.XI25.NET58_XI11.XI25.MM27_s
+ N_VDD_XI11.XI25.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=1.125e-12 AS=9.375e-13
+ PD=3e-06 PS=2.75e-06
mXI11.XI26.MM27 N_XI11.XI26.NET31_XI11.XI26.MM27_d
+ N_XI11.XI26.NET35_XI11.XI26.MM27_g N_XI11.XI26.NET58_XI11.XI26.MM27_s
+ N_VDD_XI11.XI26.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=1.125e-12 AS=9.375e-13
+ PD=3e-06 PS=2.75e-06
mXI11.XI24.MM27 N_XI11.XI24.NET31_XI11.XI24.MM27_d
+ N_XI11.XI24.NET35_XI11.XI24.MM27_g N_XI11.XI24.NET58_XI11.XI24.MM27_s
+ N_VDD_XI11.XI24.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=1.125e-12 AS=9.375e-13
+ PD=3e-06 PS=2.75e-06
mXI11.XI27.MM27 N_XI11.XI27.NET31_XI11.XI27.MM27_d
+ N_XI11.XI27.NET35_XI11.XI27.MM27_g N_XI11.XI27.NET58_XI11.XI27.MM27_s
+ N_VDD_XI11.XI27.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=1.125e-12 AS=9.375e-13
+ PD=3e-06 PS=2.75e-06
mXI11.XI22.MM27 N_XI11.XI22.NET31_XI11.XI22.MM27_d
+ N_XI11.XI22.NET35_XI11.XI22.MM27_g N_XI11.XI22.NET58_XI11.XI22.MM27_s
+ N_VDD_XI11.XI22.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=1.125e-12 AS=9.375e-13
+ PD=3e-06 PS=2.75e-06
mXI11.XI21.MM27 N_XI11.XI21.NET31_XI11.XI21.MM27_d
+ N_XI11.XI21.NET35_XI11.XI21.MM27_g N_XI11.XI21.NET58_XI11.XI21.MM27_s
+ N_VDD_XI11.XI21.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=1.125e-12 AS=9.375e-13
+ PD=3e-06 PS=2.75e-06
mXI11.XI23.MM27 N_XI11.XI23.NET31_XI11.XI23.MM27_d
+ N_XI11.XI23.NET35_XI11.XI23.MM27_g N_XI11.XI23.NET58_XI11.XI23.MM27_s
+ N_VDD_XI11.XI23.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=1.125e-12 AS=9.375e-13
+ PD=3e-06 PS=2.75e-06
mXI11.XI19.MM27 N_XI11.XI19.NET31_XI11.XI19.MM27_d
+ N_XI11.XI19.NET35_XI11.XI19.MM27_g N_XI11.XI19.NET58_XI11.XI19.MM27_s
+ N_VDD_XI11.XI19.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=1.125e-12 AS=9.375e-13
+ PD=3e-06 PS=2.75e-06
mXI11.XI20.MM27 N_XI11.XI20.NET31_XI11.XI20.MM27_d
+ N_XI11.XI20.NET35_XI11.XI20.MM27_g N_XI11.XI20.NET58_XI11.XI20.MM27_s
+ N_VDD_XI11.XI20.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=1.125e-12 AS=9.375e-13
+ PD=3e-06 PS=2.75e-06
mXI11.XI18.MM27 N_XI11.XI18.NET31_XI11.XI18.MM27_d
+ N_XI11.XI18.NET35_XI11.XI18.MM27_g N_XI11.XI18.NET58_XI11.XI18.MM27_s
+ N_VDD_XI11.XI18.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=1.125e-12 AS=9.375e-13
+ PD=3e-06 PS=2.75e-06
mXI11.XI17.MM27 N_XI11.XI17.NET31_XI11.XI17.MM27_d
+ N_XI11.XI17.NET35_XI11.XI17.MM27_g N_XI11.XI17.NET58_XI11.XI17.MM27_s
+ N_VDD_XI11.XI17.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=1.125e-12 AS=9.375e-13
+ PD=3e-06 PS=2.75e-06
mXI11.XI0.MM27 N_XI11.XI0.NET31_XI11.XI0.MM27_d N_XI11.XI0.NET35_XI11.XI0.MM27_g
+ N_XI11.XI0.NET58_XI11.XI0.MM27_s N_VDD_XI11.XI0.XI0.MM1_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.125e-12 AS=9.375e-13 PD=3e-06 PS=2.75e-06
mXI11.XI30.MM3 N_XI11.XI30.NET15_XI11.XI30.MM3_d
+ N_XI11.XI30.NET58_XI11.XI30.MM3_g N_VDD_XI11.XI30.MM3_s
+ N_VDD_XI11.XI30.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI11.XI29.MM3 N_XI11.XI29.NET15_XI11.XI29.MM3_d
+ N_XI11.XI29.NET58_XI11.XI29.MM3_g N_VDD_XI11.XI29.MM3_s
+ N_VDD_XI11.XI29.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI11.XI31.MM3 N_XI11.XI31.NET15_XI11.XI31.MM3_d
+ N_XI11.XI31.NET58_XI11.XI31.MM3_g N_VDD_XI11.XI31.MM3_s
+ N_VDD_XI11.XI31.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI11.XI28.MM3 N_XI11.XI28.NET15_XI11.XI28.MM3_d
+ N_XI11.XI28.NET58_XI11.XI28.MM3_g N_VDD_XI11.XI28.MM3_s
+ N_VDD_XI11.XI28.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI11.XI25.MM3 N_XI11.XI25.NET15_XI11.XI25.MM3_d
+ N_XI11.XI25.NET58_XI11.XI25.MM3_g N_VDD_XI11.XI25.MM3_s
+ N_VDD_XI11.XI25.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI11.XI26.MM3 N_XI11.XI26.NET15_XI11.XI26.MM3_d
+ N_XI11.XI26.NET58_XI11.XI26.MM3_g N_VDD_XI11.XI26.MM3_s
+ N_VDD_XI11.XI26.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI11.XI24.MM3 N_XI11.XI24.NET15_XI11.XI24.MM3_d
+ N_XI11.XI24.NET58_XI11.XI24.MM3_g N_VDD_XI11.XI24.MM3_s
+ N_VDD_XI11.XI24.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI11.XI27.MM3 N_XI11.XI27.NET15_XI11.XI27.MM3_d
+ N_XI11.XI27.NET58_XI11.XI27.MM3_g N_VDD_XI11.XI27.MM3_s
+ N_VDD_XI11.XI27.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI11.XI22.MM3 N_XI11.XI22.NET15_XI11.XI22.MM3_d
+ N_XI11.XI22.NET58_XI11.XI22.MM3_g N_VDD_XI11.XI22.MM3_s
+ N_VDD_XI11.XI22.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI11.XI21.MM3 N_XI11.XI21.NET15_XI11.XI21.MM3_d
+ N_XI11.XI21.NET58_XI11.XI21.MM3_g N_VDD_XI11.XI21.MM3_s
+ N_VDD_XI11.XI21.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI11.XI23.MM3 N_XI11.XI23.NET15_XI11.XI23.MM3_d
+ N_XI11.XI23.NET58_XI11.XI23.MM3_g N_VDD_XI11.XI23.MM3_s
+ N_VDD_XI11.XI23.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI11.XI19.MM3 N_XI11.XI19.NET15_XI11.XI19.MM3_d
+ N_XI11.XI19.NET58_XI11.XI19.MM3_g N_VDD_XI11.XI19.MM3_s
+ N_VDD_XI11.XI19.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI11.XI20.MM3 N_XI11.XI20.NET15_XI11.XI20.MM3_d
+ N_XI11.XI20.NET58_XI11.XI20.MM3_g N_VDD_XI11.XI20.MM3_s
+ N_VDD_XI11.XI20.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI11.XI18.MM3 N_XI11.XI18.NET15_XI11.XI18.MM3_d
+ N_XI11.XI18.NET58_XI11.XI18.MM3_g N_VDD_XI11.XI18.MM3_s
+ N_VDD_XI11.XI18.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI11.XI17.MM3 N_XI11.XI17.NET15_XI11.XI17.MM3_d
+ N_XI11.XI17.NET58_XI11.XI17.MM3_g N_VDD_XI11.XI17.MM3_s
+ N_VDD_XI11.XI17.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI11.XI0.MM3 N_XI11.XI0.NET15_XI11.XI0.MM3_d N_XI11.XI0.NET58_XI11.XI0.MM3_g
+ N_VDD_XI11.XI0.MM3_s N_VDD_XI11.XI0.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI11.XI30.MM1 N_XI11.XI30.NET54_XI11.XI30.MM1_d
+ N_XI11.XI30.NET15_XI11.XI30.MM1_g N_VDD_XI11.XI30.MM1_s
+ N_VDD_XI11.XI30.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI11.XI29.MM1 N_XI11.XI29.NET54_XI11.XI29.MM1_d
+ N_XI11.XI29.NET15_XI11.XI29.MM1_g N_VDD_XI11.XI29.MM1_s
+ N_VDD_XI11.XI29.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI11.XI31.MM1 N_XI11.XI31.NET54_XI11.XI31.MM1_d
+ N_XI11.XI31.NET15_XI11.XI31.MM1_g N_VDD_XI11.XI31.MM1_s
+ N_VDD_XI11.XI31.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI11.XI28.MM1 N_XI11.XI28.NET54_XI11.XI28.MM1_d
+ N_XI11.XI28.NET15_XI11.XI28.MM1_g N_VDD_XI11.XI28.MM1_s
+ N_VDD_XI11.XI28.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI11.XI25.MM1 N_XI11.XI25.NET54_XI11.XI25.MM1_d
+ N_XI11.XI25.NET15_XI11.XI25.MM1_g N_VDD_XI11.XI25.MM1_s
+ N_VDD_XI11.XI25.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI11.XI26.MM1 N_XI11.XI26.NET54_XI11.XI26.MM1_d
+ N_XI11.XI26.NET15_XI11.XI26.MM1_g N_VDD_XI11.XI26.MM1_s
+ N_VDD_XI11.XI26.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI11.XI24.MM1 N_XI11.XI24.NET54_XI11.XI24.MM1_d
+ N_XI11.XI24.NET15_XI11.XI24.MM1_g N_VDD_XI11.XI24.MM1_s
+ N_VDD_XI11.XI24.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI11.XI27.MM1 N_XI11.XI27.NET54_XI11.XI27.MM1_d
+ N_XI11.XI27.NET15_XI11.XI27.MM1_g N_VDD_XI11.XI27.MM1_s
+ N_VDD_XI11.XI27.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI11.XI22.MM1 N_XI11.XI22.NET54_XI11.XI22.MM1_d
+ N_XI11.XI22.NET15_XI11.XI22.MM1_g N_VDD_XI11.XI22.MM1_s
+ N_VDD_XI11.XI22.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI11.XI21.MM1 N_XI11.XI21.NET54_XI11.XI21.MM1_d
+ N_XI11.XI21.NET15_XI11.XI21.MM1_g N_VDD_XI11.XI21.MM1_s
+ N_VDD_XI11.XI21.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI11.XI23.MM1 N_XI11.XI23.NET54_XI11.XI23.MM1_d
+ N_XI11.XI23.NET15_XI11.XI23.MM1_g N_VDD_XI11.XI23.MM1_s
+ N_VDD_XI11.XI23.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI11.XI19.MM1 N_XI11.XI19.NET54_XI11.XI19.MM1_d
+ N_XI11.XI19.NET15_XI11.XI19.MM1_g N_VDD_XI11.XI19.MM1_s
+ N_VDD_XI11.XI19.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI11.XI20.MM1 N_XI11.XI20.NET54_XI11.XI20.MM1_d
+ N_XI11.XI20.NET15_XI11.XI20.MM1_g N_VDD_XI11.XI20.MM1_s
+ N_VDD_XI11.XI20.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI11.XI18.MM1 N_XI11.XI18.NET54_XI11.XI18.MM1_d
+ N_XI11.XI18.NET15_XI11.XI18.MM1_g N_VDD_XI11.XI18.MM1_s
+ N_VDD_XI11.XI18.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI11.XI17.MM1 N_XI11.XI17.NET54_XI11.XI17.MM1_d
+ N_XI11.XI17.NET15_XI11.XI17.MM1_g N_VDD_XI11.XI17.MM1_s
+ N_VDD_XI11.XI17.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI11.XI0.MM1 N_XI11.XI0.NET54_XI11.XI0.MM1_d N_XI11.XI0.NET15_XI11.XI0.MM1_g
+ N_VDD_XI11.XI0.MM1_s N_VDD_XI11.XI0.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI11.XI30.MM35 N_XI11.XI30.NET58_XI11.XI30.MM35_d
+ N_XI11.XI30.CLKB_XI11.XI30.MM35_g N_XI11.XI30.NET54_XI11.XI30.MM35_s
+ N_VDD_XI11.XI30.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI11.XI29.MM35 N_XI11.XI29.NET58_XI11.XI29.MM35_d
+ N_XI11.XI29.CLKB_XI11.XI29.MM35_g N_XI11.XI29.NET54_XI11.XI29.MM35_s
+ N_VDD_XI11.XI29.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI11.XI31.MM35 N_XI11.XI31.NET58_XI11.XI31.MM35_d
+ N_XI11.XI31.CLKB_XI11.XI31.MM35_g N_XI11.XI31.NET54_XI11.XI31.MM35_s
+ N_VDD_XI11.XI31.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI11.XI28.MM35 N_XI11.XI28.NET58_XI11.XI28.MM35_d
+ N_XI11.XI28.CLKB_XI11.XI28.MM35_g N_XI11.XI28.NET54_XI11.XI28.MM35_s
+ N_VDD_XI11.XI28.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI11.XI25.MM35 N_XI11.XI25.NET58_XI11.XI25.MM35_d
+ N_XI11.XI25.CLKB_XI11.XI25.MM35_g N_XI11.XI25.NET54_XI11.XI25.MM35_s
+ N_VDD_XI11.XI25.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI11.XI26.MM35 N_XI11.XI26.NET58_XI11.XI26.MM35_d
+ N_XI11.XI26.CLKB_XI11.XI26.MM35_g N_XI11.XI26.NET54_XI11.XI26.MM35_s
+ N_VDD_XI11.XI26.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI11.XI24.MM35 N_XI11.XI24.NET58_XI11.XI24.MM35_d
+ N_XI11.XI24.CLKB_XI11.XI24.MM35_g N_XI11.XI24.NET54_XI11.XI24.MM35_s
+ N_VDD_XI11.XI24.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI11.XI27.MM35 N_XI11.XI27.NET58_XI11.XI27.MM35_d
+ N_XI11.XI27.CLKB_XI11.XI27.MM35_g N_XI11.XI27.NET54_XI11.XI27.MM35_s
+ N_VDD_XI11.XI27.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI11.XI22.MM35 N_XI11.XI22.NET58_XI11.XI22.MM35_d
+ N_XI11.XI22.CLKB_XI11.XI22.MM35_g N_XI11.XI22.NET54_XI11.XI22.MM35_s
+ N_VDD_XI11.XI22.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI11.XI21.MM35 N_XI11.XI21.NET58_XI11.XI21.MM35_d
+ N_XI11.XI21.CLKB_XI11.XI21.MM35_g N_XI11.XI21.NET54_XI11.XI21.MM35_s
+ N_VDD_XI11.XI21.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI11.XI23.MM35 N_XI11.XI23.NET58_XI11.XI23.MM35_d
+ N_XI11.XI23.CLKB_XI11.XI23.MM35_g N_XI11.XI23.NET54_XI11.XI23.MM35_s
+ N_VDD_XI11.XI23.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI11.XI19.MM35 N_XI11.XI19.NET58_XI11.XI19.MM35_d
+ N_XI11.XI19.CLKB_XI11.XI19.MM35_g N_XI11.XI19.NET54_XI11.XI19.MM35_s
+ N_VDD_XI11.XI19.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI11.XI20.MM35 N_XI11.XI20.NET58_XI11.XI20.MM35_d
+ N_XI11.XI20.CLKB_XI11.XI20.MM35_g N_XI11.XI20.NET54_XI11.XI20.MM35_s
+ N_VDD_XI11.XI20.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI11.XI18.MM35 N_XI11.XI18.NET58_XI11.XI18.MM35_d
+ N_XI11.XI18.CLKB_XI11.XI18.MM35_g N_XI11.XI18.NET54_XI11.XI18.MM35_s
+ N_VDD_XI11.XI18.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI11.XI17.MM35 N_XI11.XI17.NET58_XI11.XI17.MM35_d
+ N_XI11.XI17.CLKB_XI11.XI17.MM35_g N_XI11.XI17.NET54_XI11.XI17.MM35_s
+ N_VDD_XI11.XI17.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI11.XI0.MM35 N_XI11.XI0.NET58_XI11.XI0.MM35_d N_XI11.XI0.CLKB_XI11.XI0.MM35_g
+ N_XI11.XI0.NET54_XI11.XI0.MM35_s N_VDD_XI11.XI0.XI0.MM1_b P_18 L=1.8e-07
+ W=1.5e-06 AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI11.XI30.MM37 N_XI11.XI30.NET15_XI11.XI30.MM37_d
+ N_XI11.XI30.CLKB_XI11.XI30.MM37_g N_XI11.XI30.NET14_XI11.XI30.MM37_s
+ N_VDD_XI11.XI30.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=1.125e-12 AS=9.375e-13
+ PD=3e-06 PS=2.75e-06
mXI11.XI29.MM37 N_XI11.XI29.NET15_XI11.XI29.MM37_d
+ N_XI11.XI29.CLKB_XI11.XI29.MM37_g N_XI11.XI29.NET14_XI11.XI29.MM37_s
+ N_VDD_XI11.XI29.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=1.125e-12 AS=9.375e-13
+ PD=3e-06 PS=2.75e-06
mXI11.XI31.MM37 N_XI11.XI31.NET15_XI11.XI31.MM37_d
+ N_XI11.XI31.CLKB_XI11.XI31.MM37_g N_XI11.XI31.NET14_XI11.XI31.MM37_s
+ N_VDD_XI11.XI31.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=1.125e-12 AS=9.375e-13
+ PD=3e-06 PS=2.75e-06
mXI11.XI28.MM37 N_XI11.XI28.NET15_XI11.XI28.MM37_d
+ N_XI11.XI28.CLKB_XI11.XI28.MM37_g N_XI11.XI28.NET14_XI11.XI28.MM37_s
+ N_VDD_XI11.XI28.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=1.125e-12 AS=9.375e-13
+ PD=3e-06 PS=2.75e-06
mXI11.XI25.MM37 N_XI11.XI25.NET15_XI11.XI25.MM37_d
+ N_XI11.XI25.CLKB_XI11.XI25.MM37_g N_XI11.XI25.NET14_XI11.XI25.MM37_s
+ N_VDD_XI11.XI25.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=1.125e-12 AS=9.375e-13
+ PD=3e-06 PS=2.75e-06
mXI11.XI26.MM37 N_XI11.XI26.NET15_XI11.XI26.MM37_d
+ N_XI11.XI26.CLKB_XI11.XI26.MM37_g N_XI11.XI26.NET14_XI11.XI26.MM37_s
+ N_VDD_XI11.XI26.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=1.125e-12 AS=9.375e-13
+ PD=3e-06 PS=2.75e-06
mXI11.XI24.MM37 N_XI11.XI24.NET15_XI11.XI24.MM37_d
+ N_XI11.XI24.CLKB_XI11.XI24.MM37_g N_XI11.XI24.NET14_XI11.XI24.MM37_s
+ N_VDD_XI11.XI24.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=1.125e-12 AS=9.375e-13
+ PD=3e-06 PS=2.75e-06
mXI11.XI27.MM37 N_XI11.XI27.NET15_XI11.XI27.MM37_d
+ N_XI11.XI27.CLKB_XI11.XI27.MM37_g N_XI11.XI27.NET14_XI11.XI27.MM37_s
+ N_VDD_XI11.XI27.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=1.125e-12 AS=9.375e-13
+ PD=3e-06 PS=2.75e-06
mXI11.XI22.MM37 N_XI11.XI22.NET15_XI11.XI22.MM37_d
+ N_XI11.XI22.CLKB_XI11.XI22.MM37_g N_XI11.XI22.NET14_XI11.XI22.MM37_s
+ N_VDD_XI11.XI22.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=1.125e-12 AS=9.375e-13
+ PD=3e-06 PS=2.75e-06
mXI11.XI21.MM37 N_XI11.XI21.NET15_XI11.XI21.MM37_d
+ N_XI11.XI21.CLKB_XI11.XI21.MM37_g N_XI11.XI21.NET14_XI11.XI21.MM37_s
+ N_VDD_XI11.XI21.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=1.125e-12 AS=9.375e-13
+ PD=3e-06 PS=2.75e-06
mXI11.XI23.MM37 N_XI11.XI23.NET15_XI11.XI23.MM37_d
+ N_XI11.XI23.CLKB_XI11.XI23.MM37_g N_XI11.XI23.NET14_XI11.XI23.MM37_s
+ N_VDD_XI11.XI23.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=1.125e-12 AS=9.375e-13
+ PD=3e-06 PS=2.75e-06
mXI11.XI19.MM37 N_XI11.XI19.NET15_XI11.XI19.MM37_d
+ N_XI11.XI19.CLKB_XI11.XI19.MM37_g N_XI11.XI19.NET14_XI11.XI19.MM37_s
+ N_VDD_XI11.XI19.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=1.125e-12 AS=9.375e-13
+ PD=3e-06 PS=2.75e-06
mXI11.XI20.MM37 N_XI11.XI20.NET15_XI11.XI20.MM37_d
+ N_XI11.XI20.CLKB_XI11.XI20.MM37_g N_XI11.XI20.NET14_XI11.XI20.MM37_s
+ N_VDD_XI11.XI20.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=1.125e-12 AS=9.375e-13
+ PD=3e-06 PS=2.75e-06
mXI11.XI18.MM37 N_XI11.XI18.NET15_XI11.XI18.MM37_d
+ N_XI11.XI18.CLKB_XI11.XI18.MM37_g N_XI11.XI18.NET14_XI11.XI18.MM37_s
+ N_VDD_XI11.XI18.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=1.125e-12 AS=9.375e-13
+ PD=3e-06 PS=2.75e-06
mXI11.XI17.MM37 N_XI11.XI17.NET15_XI11.XI17.MM37_d
+ N_XI11.XI17.CLKB_XI11.XI17.MM37_g N_XI11.XI17.NET14_XI11.XI17.MM37_s
+ N_VDD_XI11.XI17.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=1.125e-12 AS=9.375e-13
+ PD=3e-06 PS=2.75e-06
mXI11.XI0.MM37 N_XI11.XI0.NET15_XI11.XI0.MM37_d N_XI11.XI0.CLKB_XI11.XI0.MM37_g
+ N_XI11.XI0.NET14_XI11.XI0.MM37_s N_VDD_XI11.XI0.XI0.MM1_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.125e-12 AS=9.375e-13 PD=3e-06 PS=2.75e-06
mXI11.XI30.MM13 N_ACC15_XI11.XI30.MM13_d N_XI11.XI30.NET14_XI11.XI30.MM13_g
+ N_VDD_XI11.XI30.MM13_s N_VDD_XI11.XI30.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI11.XI29.MM13 N_ACC14_XI11.XI29.MM13_d N_XI11.XI29.NET14_XI11.XI29.MM13_g
+ N_VDD_XI11.XI29.MM13_s N_VDD_XI11.XI29.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI11.XI31.MM13 N_ACC13_XI11.XI31.MM13_d N_XI11.XI31.NET14_XI11.XI31.MM13_g
+ N_VDD_XI11.XI31.MM13_s N_VDD_XI11.XI31.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI11.XI28.MM13 N_ACC12_XI11.XI28.MM13_d N_XI11.XI28.NET14_XI11.XI28.MM13_g
+ N_VDD_XI11.XI28.MM13_s N_VDD_XI11.XI28.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI11.XI25.MM13 N_ACC11_XI11.XI25.MM13_d N_XI11.XI25.NET14_XI11.XI25.MM13_g
+ N_VDD_XI11.XI25.MM13_s N_VDD_XI11.XI25.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI11.XI26.MM13 N_ACC10_XI11.XI26.MM13_d N_XI11.XI26.NET14_XI11.XI26.MM13_g
+ N_VDD_XI11.XI26.MM13_s N_VDD_XI11.XI26.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI11.XI24.MM13 N_ACC9_XI11.XI24.MM13_d N_XI11.XI24.NET14_XI11.XI24.MM13_g
+ N_VDD_XI11.XI24.MM13_s N_VDD_XI11.XI24.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI11.XI27.MM13 N_ACC8_XI11.XI27.MM13_d N_XI11.XI27.NET14_XI11.XI27.MM13_g
+ N_VDD_XI11.XI27.MM13_s N_VDD_XI11.XI27.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI11.XI22.MM13 N_ACC7_XI11.XI22.MM13_d N_XI11.XI22.NET14_XI11.XI22.MM13_g
+ N_VDD_XI11.XI22.MM13_s N_VDD_XI11.XI22.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI11.XI21.MM13 N_ACC6_XI11.XI21.MM13_d N_XI11.XI21.NET14_XI11.XI21.MM13_g
+ N_VDD_XI11.XI21.MM13_s N_VDD_XI11.XI21.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI11.XI23.MM13 N_ACC5_XI11.XI23.MM13_d N_XI11.XI23.NET14_XI11.XI23.MM13_g
+ N_VDD_XI11.XI23.MM13_s N_VDD_XI11.XI23.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI11.XI19.MM13 N_ACC4_XI11.XI19.MM13_d N_XI11.XI19.NET14_XI11.XI19.MM13_g
+ N_VDD_XI11.XI19.MM13_s N_VDD_XI11.XI19.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI11.XI20.MM13 N_ACC3_XI11.XI20.MM13_d N_XI11.XI20.NET14_XI11.XI20.MM13_g
+ N_VDD_XI11.XI20.MM13_s N_VDD_XI11.XI20.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI11.XI18.MM13 N_ACC2_XI11.XI18.MM13_d N_XI11.XI18.NET14_XI11.XI18.MM13_g
+ N_VDD_XI11.XI18.MM13_s N_VDD_XI11.XI18.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI11.XI17.MM13 N_ACC1_XI11.XI17.MM13_d N_XI11.XI17.NET14_XI11.XI17.MM13_g
+ N_VDD_XI11.XI17.MM13_s N_VDD_XI11.XI17.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI11.XI0.MM13 N_ACC0_XI11.XI0.MM13_d N_XI11.XI0.NET14_XI11.XI0.MM13_g
+ N_VDD_XI11.XI0.MM13_s N_VDD_XI11.XI0.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI11.XI30.MM14 N_XI11.BAR_Q16_XI11.XI30.MM14_d N_ACC15_XI11.XI30.MM14_g
+ N_VDD_XI11.XI30.MM14_s N_VDD_XI11.XI30.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI11.XI29.MM14 N_XI11.BAR_Q15_XI11.XI29.MM14_d N_ACC14_XI11.XI29.MM14_g
+ N_VDD_XI11.XI29.MM14_s N_VDD_XI11.XI29.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI11.XI31.MM14 N_XI11.BAR_Q14_XI11.XI31.MM14_d N_ACC13_XI11.XI31.MM14_g
+ N_VDD_XI11.XI31.MM14_s N_VDD_XI11.XI31.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI11.XI28.MM14 N_XI11.BAR_Q13_XI11.XI28.MM14_d N_ACC12_XI11.XI28.MM14_g
+ N_VDD_XI11.XI28.MM14_s N_VDD_XI11.XI28.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI11.XI25.MM14 N_XI11.BAR_Q12_XI11.XI25.MM14_d N_ACC11_XI11.XI25.MM14_g
+ N_VDD_XI11.XI25.MM14_s N_VDD_XI11.XI25.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI11.XI26.MM14 N_XI11.BAR_Q11_XI11.XI26.MM14_d N_ACC10_XI11.XI26.MM14_g
+ N_VDD_XI11.XI26.MM14_s N_VDD_XI11.XI26.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI11.XI24.MM14 N_XI11.BAR_Q10_XI11.XI24.MM14_d N_ACC9_XI11.XI24.MM14_g
+ N_VDD_XI11.XI24.MM14_s N_VDD_XI11.XI24.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI11.XI27.MM14 N_XI11.BAR_Q9_XI11.XI27.MM14_d N_ACC8_XI11.XI27.MM14_g
+ N_VDD_XI11.XI27.MM14_s N_VDD_XI11.XI27.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI11.XI22.MM14 N_XI11.BAR_Q8_XI11.XI22.MM14_d N_ACC7_XI11.XI22.MM14_g
+ N_VDD_XI11.XI22.MM14_s N_VDD_XI11.XI22.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI11.XI21.MM14 N_XI11.BAR_Q7_XI11.XI21.MM14_d N_ACC6_XI11.XI21.MM14_g
+ N_VDD_XI11.XI21.MM14_s N_VDD_XI11.XI21.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI11.XI23.MM14 N_XI11.BAR_Q6_XI11.XI23.MM14_d N_ACC5_XI11.XI23.MM14_g
+ N_VDD_XI11.XI23.MM14_s N_VDD_XI11.XI23.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI11.XI19.MM14 N_XI11.BAR_Q5_XI11.XI19.MM14_d N_ACC4_XI11.XI19.MM14_g
+ N_VDD_XI11.XI19.MM14_s N_VDD_XI11.XI19.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI11.XI20.MM14 N_XI11.BAR_Q4_XI11.XI20.MM14_d N_ACC3_XI11.XI20.MM14_g
+ N_VDD_XI11.XI20.MM14_s N_VDD_XI11.XI20.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI11.XI18.MM14 N_XI11.BAR_Q3_XI11.XI18.MM14_d N_ACC2_XI11.XI18.MM14_g
+ N_VDD_XI11.XI18.MM14_s N_VDD_XI11.XI18.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI11.XI17.MM14 N_XI11.BAR_Q2_XI11.XI17.MM14_d N_ACC1_XI11.XI17.MM14_g
+ N_VDD_XI11.XI17.MM14_s N_VDD_XI11.XI17.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI11.XI0.MM14 N_XI11.BAR_Q1_XI11.XI0.MM14_d N_ACC0_XI11.XI0.MM14_g
+ N_VDD_XI11.XI0.MM14_s N_VDD_XI11.XI0.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI11.XI30.MM39 N_XI11.XI30.NET14_XI11.XI30.MM39_d
+ N_XI11.XI30.NET35_XI11.XI30.MM39_g N_XI11.BAR_Q16_XI11.XI30.MM39_s
+ N_VDD_XI11.XI30.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI11.XI29.MM39 N_XI11.XI29.NET14_XI11.XI29.MM39_d
+ N_XI11.XI29.NET35_XI11.XI29.MM39_g N_XI11.BAR_Q15_XI11.XI29.MM39_s
+ N_VDD_XI11.XI29.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI11.XI31.MM39 N_XI11.XI31.NET14_XI11.XI31.MM39_d
+ N_XI11.XI31.NET35_XI11.XI31.MM39_g N_XI11.BAR_Q14_XI11.XI31.MM39_s
+ N_VDD_XI11.XI31.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI11.XI28.MM39 N_XI11.XI28.NET14_XI11.XI28.MM39_d
+ N_XI11.XI28.NET35_XI11.XI28.MM39_g N_XI11.BAR_Q13_XI11.XI28.MM39_s
+ N_VDD_XI11.XI28.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI11.XI25.MM39 N_XI11.XI25.NET14_XI11.XI25.MM39_d
+ N_XI11.XI25.NET35_XI11.XI25.MM39_g N_XI11.BAR_Q12_XI11.XI25.MM39_s
+ N_VDD_XI11.XI25.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI11.XI26.MM39 N_XI11.XI26.NET14_XI11.XI26.MM39_d
+ N_XI11.XI26.NET35_XI11.XI26.MM39_g N_XI11.BAR_Q11_XI11.XI26.MM39_s
+ N_VDD_XI11.XI26.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI11.XI24.MM39 N_XI11.XI24.NET14_XI11.XI24.MM39_d
+ N_XI11.XI24.NET35_XI11.XI24.MM39_g N_XI11.BAR_Q10_XI11.XI24.MM39_s
+ N_VDD_XI11.XI24.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI11.XI27.MM39 N_XI11.XI27.NET14_XI11.XI27.MM39_d
+ N_XI11.XI27.NET35_XI11.XI27.MM39_g N_XI11.BAR_Q9_XI11.XI27.MM39_s
+ N_VDD_XI11.XI27.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI11.XI22.MM39 N_XI11.XI22.NET14_XI11.XI22.MM39_d
+ N_XI11.XI22.NET35_XI11.XI22.MM39_g N_XI11.BAR_Q8_XI11.XI22.MM39_s
+ N_VDD_XI11.XI22.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI11.XI21.MM39 N_XI11.XI21.NET14_XI11.XI21.MM39_d
+ N_XI11.XI21.NET35_XI11.XI21.MM39_g N_XI11.BAR_Q7_XI11.XI21.MM39_s
+ N_VDD_XI11.XI21.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI11.XI23.MM39 N_XI11.XI23.NET14_XI11.XI23.MM39_d
+ N_XI11.XI23.NET35_XI11.XI23.MM39_g N_XI11.BAR_Q6_XI11.XI23.MM39_s
+ N_VDD_XI11.XI23.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI11.XI19.MM39 N_XI11.XI19.NET14_XI11.XI19.MM39_d
+ N_XI11.XI19.NET35_XI11.XI19.MM39_g N_XI11.BAR_Q5_XI11.XI19.MM39_s
+ N_VDD_XI11.XI19.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI11.XI20.MM39 N_XI11.XI20.NET14_XI11.XI20.MM39_d
+ N_XI11.XI20.NET35_XI11.XI20.MM39_g N_XI11.BAR_Q4_XI11.XI20.MM39_s
+ N_VDD_XI11.XI20.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI11.XI18.MM39 N_XI11.XI18.NET14_XI11.XI18.MM39_d
+ N_XI11.XI18.NET35_XI11.XI18.MM39_g N_XI11.BAR_Q3_XI11.XI18.MM39_s
+ N_VDD_XI11.XI18.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI11.XI17.MM39 N_XI11.XI17.NET14_XI11.XI17.MM39_d
+ N_XI11.XI17.NET35_XI11.XI17.MM39_g N_XI11.BAR_Q2_XI11.XI17.MM39_s
+ N_VDD_XI11.XI17.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI11.XI0.MM39 N_XI11.XI0.NET14_XI11.XI0.MM39_d N_XI11.XI0.NET35_XI11.XI0.MM39_g
+ N_XI11.BAR_Q1_XI11.XI0.MM39_s N_VDD_XI11.XI0.XI0.MM1_b P_18 L=1.8e-07
+ W=1.5e-06 AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI20.XI11.MM1 N_NET594_XI20.XI11.MM1_d N_NET241_XI20.XI11.MM1_g
+ N_VDD_XI20.XI11.MM1_s N_VDD_XI20.XI11.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI21.XI11.MM1 N_NET628_XI21.XI11.MM1_d N_NET241_XI21.XI11.MM1_g
+ N_VDD_XI21.XI11.MM1_s N_VDD_XI20.XI11.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI20.XI12.MM1 N_NET595_XI20.XI12.MM1_d N_NET242_XI20.XI12.MM1_g
+ N_VDD_XI20.XI12.MM1_s N_VDD_XI20.XI11.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI21.XI12.MM1 N_NET629_XI21.XI12.MM1_d N_NET242_XI21.XI12.MM1_g
+ N_VDD_XI21.XI12.MM1_s N_VDD_XI20.XI11.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI20.XI10.MM1 N_NET596_XI20.XI10.MM1_d N_NET243_XI20.XI10.MM1_g
+ N_VDD_XI20.XI10.MM1_s N_VDD_XI20.XI11.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI21.XI10.MM1 N_NET630_XI21.XI10.MM1_d N_NET243_XI21.XI10.MM1_g
+ N_VDD_XI21.XI10.MM1_s N_VDD_XI20.XI11.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI20.XI9.MM1 N_NET597_XI20.XI9.MM1_d N_NET244_XI20.XI9.MM1_g
+ N_VDD_XI20.XI9.MM1_s N_VDD_XI20.XI11.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI21.XI9.MM1 N_NET631_XI21.XI9.MM1_d N_NET244_XI21.XI9.MM1_g
+ N_VDD_XI21.XI9.MM1_s N_VDD_XI20.XI11.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI20.XI14.MM1 N_NET598_XI20.XI14.MM1_d N_NET245_XI20.XI14.MM1_g
+ N_VDD_XI20.XI14.MM1_s N_VDD_XI20.XI11.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI21.XI14.MM1 N_NET632_XI21.XI14.MM1_d N_NET245_XI21.XI14.MM1_g
+ N_VDD_XI21.XI14.MM1_s N_VDD_XI20.XI11.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI20.XI13.MM1 N_NET599_XI20.XI13.MM1_d N_NET246_XI20.XI13.MM1_g
+ N_VDD_XI20.XI13.MM1_s N_VDD_XI20.XI11.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI21.XI13.MM1 N_NET633_XI21.XI13.MM1_d N_NET246_XI21.XI13.MM1_g
+ N_VDD_XI21.XI13.MM1_s N_VDD_XI20.XI11.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI20.XI15.MM1 N_NET600_XI20.XI15.MM1_d N_NET247_XI20.XI15.MM1_g
+ N_VDD_XI20.XI15.MM1_s N_VDD_XI20.XI11.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI21.XI15.MM1 N_NET634_XI21.XI15.MM1_d N_NET247_XI21.XI15.MM1_g
+ N_VDD_XI21.XI15.MM1_s N_VDD_XI20.XI11.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI20.XI6.MM1 N_NET601_XI20.XI6.MM1_d N_NET248_XI20.XI6.MM1_g
+ N_VDD_XI20.XI6.MM1_s N_VDD_XI20.XI11.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI21.XI6.MM1 N_NET635_XI21.XI6.MM1_d N_NET248_XI21.XI6.MM1_g
+ N_VDD_XI21.XI6.MM1_s N_VDD_XI20.XI11.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI20.XI5.MM1 N_NET602_XI20.XI5.MM1_d N_NET249_XI20.XI5.MM1_g
+ N_VDD_XI20.XI5.MM1_s N_VDD_XI20.XI11.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI21.XI5.MM1 N_NET636_XI21.XI5.MM1_d N_NET249_XI21.XI5.MM1_g
+ N_VDD_XI21.XI5.MM1_s N_VDD_XI20.XI11.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI20.XI7.MM1 N_NET603_XI20.XI7.MM1_d N_NET250_XI20.XI7.MM1_g
+ N_VDD_XI20.XI7.MM1_s N_VDD_XI20.XI11.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI21.XI7.MM1 N_NET637_XI21.XI7.MM1_d N_NET250_XI21.XI7.MM1_g
+ N_VDD_XI21.XI7.MM1_s N_VDD_XI20.XI11.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI20.XI8.MM1 N_NET604_XI20.XI8.MM1_d N_NET251_XI20.XI8.MM1_g
+ N_VDD_XI20.XI8.MM1_s N_VDD_XI20.XI11.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI21.XI8.MM1 N_NET638_XI21.XI8.MM1_d N_NET251_XI21.XI8.MM1_g
+ N_VDD_XI21.XI8.MM1_s N_VDD_XI20.XI11.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI20.XI3.MM1 N_NET605_XI20.XI3.MM1_d N_NET252_XI20.XI3.MM1_g
+ N_VDD_XI20.XI3.MM1_s N_VDD_XI20.XI11.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI21.XI3.MM1 N_NET639_XI21.XI3.MM1_d N_NET252_XI21.XI3.MM1_g
+ N_VDD_XI21.XI3.MM1_s N_VDD_XI20.XI11.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI20.XI4.MM1 N_NET606_XI20.XI4.MM1_d N_NET253_XI20.XI4.MM1_g
+ N_VDD_XI20.XI4.MM1_s N_VDD_XI20.XI11.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI21.XI4.MM1 N_NET640_XI21.XI4.MM1_d N_NET253_XI21.XI4.MM1_g
+ N_VDD_XI21.XI4.MM1_s N_VDD_XI20.XI11.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI20.XI2.MM1 N_NET607_XI20.XI2.MM1_d N_NET254_XI20.XI2.MM1_g
+ N_VDD_XI20.XI2.MM1_s N_VDD_XI20.XI11.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI21.XI2.MM1 N_NET641_XI21.XI2.MM1_d N_NET254_XI21.XI2.MM1_g
+ N_VDD_XI21.XI2.MM1_s N_VDD_XI20.XI11.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI20.XI1.MM1 N_NET608_XI20.XI1.MM1_d N_NET255_XI20.XI1.MM1_g
+ N_VDD_XI20.XI1.MM1_s N_VDD_XI20.XI11.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI21.XI1.MM1 N_NET642_XI21.XI1.MM1_d N_NET255_XI21.XI1.MM1_g
+ N_VDD_XI21.XI1.MM1_s N_VDD_XI20.XI11.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI20.XI0.MM1 N_NET609_XI20.XI0.MM1_d N_NET256_XI20.XI0.MM1_g
+ N_VDD_XI20.XI0.MM1_s N_VDD_XI20.XI11.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI21.XI0.MM1 N_NET643_XI21.XI0.MM1_d N_NET256_XI21.XI0.MM1_g
+ N_VDD_XI21.XI0.MM1_s N_VDD_XI20.XI11.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI0.XI134.XI9.MM1 N_XI0.XI134.NET43_XI0.XI134.XI9.MM1_d
+ N_NET594_XI0.XI134.XI9.MM1_g N_VDD_XI0.XI134.XI9.MM1_s
+ N_VDD_XI0.XI134.XI9.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI0.XI153.XI1.MM3 N_XI0.XI153.NET6_XI0.XI153.XI1.MM3_d
+ N_NET595_XI0.XI153.XI1.MM3_g N_VDD_XI0.XI153.XI1.MM3_s
+ N_VDD_XI0.XI153.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.35e-13
+ PD=7.4e-07 PS=2.48e-06
mXI0.XI154.XI1.MM3 N_XI0.XI154.NET6_XI0.XI154.XI1.MM3_d
+ N_NET596_XI0.XI154.XI1.MM3_g N_VDD_XI0.XI154.XI1.MM3_s
+ N_VDD_XI0.XI154.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.35e-13
+ PD=7.4e-07 PS=2.48e-06
mXI0.XI157.XI1.MM3 N_XI0.XI157.NET6_XI0.XI157.XI1.MM3_d
+ N_NET597_XI0.XI157.XI1.MM3_g N_VDD_XI0.XI157.XI1.MM3_s
+ N_VDD_XI0.XI157.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.35e-13
+ PD=7.4e-07 PS=2.48e-06
mXI0.XI156.XI1.MM3 N_XI0.XI156.NET6_XI0.XI156.XI1.MM3_d
+ N_NET598_XI0.XI156.XI1.MM3_g N_VDD_XI0.XI156.XI1.MM3_s
+ N_VDD_XI0.XI156.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.35e-13
+ PD=7.4e-07 PS=2.48e-06
mXI0.XI155.XI1.MM3 N_XI0.XI155.NET6_XI0.XI155.XI1.MM3_d
+ N_NET599_XI0.XI155.XI1.MM3_g N_VDD_XI0.XI155.XI1.MM3_s
+ N_VDD_XI0.XI155.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.35e-13
+ PD=7.4e-07 PS=2.48e-06
mXI0.XI133.XI1.MM3 N_XI0.XI133.NET6_XI0.XI133.XI1.MM3_d
+ N_NET600_XI0.XI133.XI1.MM3_g N_VDD_XI0.XI133.XI1.MM3_s
+ N_VDD_XI0.XI133.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.35e-13
+ PD=7.4e-07 PS=2.48e-06
mXI0.XI132.XI1.MM3 N_XI0.XI132.NET6_XI0.XI132.XI1.MM3_d
+ N_NET601_XI0.XI132.XI1.MM3_g N_VDD_XI0.XI132.XI1.MM3_s
+ N_VDD_XI0.XI132.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.35e-13
+ PD=7.4e-07 PS=2.48e-06
mXI0.XI131.XI1.MM3 N_XI0.XI131.NET6_XI0.XI131.XI1.MM3_d
+ N_NET602_XI0.XI131.XI1.MM3_g N_VDD_XI0.XI131.XI1.MM3_s
+ N_VDD_XI0.XI131.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.35e-13
+ PD=7.4e-07 PS=2.48e-06
mXI0.XI111.XI1.MM3 N_XI0.XI111.NET6_XI0.XI111.XI1.MM3_d
+ N_NET603_XI0.XI111.XI1.MM3_g N_VDD_XI0.XI111.XI1.MM3_s
+ N_VDD_XI0.XI111.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.35e-13
+ PD=7.4e-07 PS=2.48e-06
mXI0.XI110.XI1.MM3 N_XI0.XI110.NET6_XI0.XI110.XI1.MM3_d
+ N_NET604_XI0.XI110.XI1.MM3_g N_VDD_XI0.XI110.XI1.MM3_s
+ N_VDD_XI0.XI110.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.35e-13
+ PD=7.4e-07 PS=2.48e-06
mXI0.XI103.XI1.MM3 N_XI0.XI103.NET6_XI0.XI103.XI1.MM3_d
+ N_NET605_XI0.XI103.XI1.MM3_g N_VDD_XI0.XI103.XI1.MM3_s
+ N_VDD_XI0.XI103.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.35e-13
+ PD=7.4e-07 PS=2.48e-06
mXI0.XI102.XI1.MM3 N_XI0.XI102.NET6_XI0.XI102.XI1.MM3_d
+ N_NET606_XI0.XI102.XI1.MM3_g N_VDD_XI0.XI102.XI1.MM3_s
+ N_VDD_XI0.XI102.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.35e-13
+ PD=7.4e-07 PS=2.48e-06
mXI0.XI88.XI1.MM3 N_XI0.XI88.NET6_XI0.XI88.XI1.MM3_d N_NET607_XI0.XI88.XI1.MM3_g
+ N_VDD_XI0.XI88.XI1.MM3_s N_VDD_XI0.XI88.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=5.55e-13 AS=7.35e-13 PD=7.4e-07 PS=2.48e-06
mXI0.XI82.XI1.MM3 N_XI0.XI82.NET6_XI0.XI82.XI1.MM3_d N_NET608_XI0.XI82.XI1.MM3_g
+ N_VDD_XI0.XI82.XI1.MM3_s N_VDD_XI0.XI82.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=5.55e-13 AS=7.35e-13 PD=7.4e-07 PS=2.48e-06
mXI0.XI10.XI1.MM3 N_XI0.XI10.NET6_XI0.XI10.XI1.MM3_d N_NET609_XI0.XI10.XI1.MM3_g
+ N_VDD_XI0.XI10.XI1.MM3_s N_VDD_XI0.XI10.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=5.55e-13 AS=7.35e-13 PD=7.4e-07 PS=2.48e-06
mXI6.MM1 N_NET0859_XI6.MM1_d N_NET0858_XI6.MM1_g N_VDD_XI6.MM1_s N_VDD_XI6.MM1_b
+ P_18 L=1.8e-07 W=9e-06 AD=4.41e-12 AS=4.41e-12 PD=9.98e-06 PS=9.98e-06
mXI0.XI153.XI1.MM1 N_XI0.XI153.NET6_XI0.XI153.XI1.MM1_d
+ N_MIN14_XI0.XI153.XI1.MM1_g N_VDD_XI0.XI153.XI1.MM1_s
+ N_VDD_XI0.XI153.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.65e-13
+ PD=7.4e-07 PS=2.52e-06
mXI0.XI154.XI1.MM1 N_XI0.XI154.NET6_XI0.XI154.XI1.MM1_d
+ N_MIN13_XI0.XI154.XI1.MM1_g N_VDD_XI0.XI154.XI1.MM1_s
+ N_VDD_XI0.XI154.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.65e-13
+ PD=7.4e-07 PS=2.52e-06
mXI0.XI157.XI1.MM1 N_XI0.XI157.NET6_XI0.XI157.XI1.MM1_d
+ N_MIN12_XI0.XI157.XI1.MM1_g N_VDD_XI0.XI157.XI1.MM1_s
+ N_VDD_XI0.XI157.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.65e-13
+ PD=7.4e-07 PS=2.52e-06
mXI0.XI156.XI1.MM1 N_XI0.XI156.NET6_XI0.XI156.XI1.MM1_d
+ N_MIN11_XI0.XI156.XI1.MM1_g N_VDD_XI0.XI156.XI1.MM1_s
+ N_VDD_XI0.XI156.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.65e-13
+ PD=7.4e-07 PS=2.52e-06
mXI0.XI155.XI1.MM1 N_XI0.XI155.NET6_XI0.XI155.XI1.MM1_d
+ N_MIN10_XI0.XI155.XI1.MM1_g N_VDD_XI0.XI155.XI1.MM1_s
+ N_VDD_XI0.XI155.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.65e-13
+ PD=7.4e-07 PS=2.52e-06
mXI0.XI133.XI1.MM1 N_XI0.XI133.NET6_XI0.XI133.XI1.MM1_d
+ N_MIN9_XI0.XI133.XI1.MM1_g N_VDD_XI0.XI133.XI1.MM1_s N_VDD_XI0.XI133.XI1.MM3_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.65e-13 PD=7.4e-07 PS=2.52e-06
mXI0.XI132.XI1.MM1 N_XI0.XI132.NET6_XI0.XI132.XI1.MM1_d
+ N_MIN8_XI0.XI132.XI1.MM1_g N_VDD_XI0.XI132.XI1.MM1_s N_VDD_XI0.XI132.XI1.MM3_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.65e-13 PD=7.4e-07 PS=2.52e-06
mXI0.XI131.XI1.MM1 N_XI0.XI131.NET6_XI0.XI131.XI1.MM1_d
+ N_MIN7_XI0.XI131.XI1.MM1_g N_VDD_XI0.XI131.XI1.MM1_s N_VDD_XI0.XI131.XI1.MM3_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.65e-13 PD=7.4e-07 PS=2.52e-06
mXI0.XI111.XI1.MM1 N_XI0.XI111.NET6_XI0.XI111.XI1.MM1_d
+ N_MIN6_XI0.XI111.XI1.MM1_g N_VDD_XI0.XI111.XI1.MM1_s N_VDD_XI0.XI111.XI1.MM3_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.65e-13 PD=7.4e-07 PS=2.52e-06
mXI0.XI110.XI1.MM1 N_XI0.XI110.NET6_XI0.XI110.XI1.MM1_d
+ N_MIN5_XI0.XI110.XI1.MM1_g N_VDD_XI0.XI110.XI1.MM1_s N_VDD_XI0.XI110.XI1.MM3_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.65e-13 PD=7.4e-07 PS=2.52e-06
mXI0.XI103.XI1.MM1 N_XI0.XI103.NET6_XI0.XI103.XI1.MM1_d
+ N_MIN4_XI0.XI103.XI1.MM1_g N_VDD_XI0.XI103.XI1.MM1_s N_VDD_XI0.XI103.XI1.MM3_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.65e-13 PD=7.4e-07 PS=2.52e-06
mXI0.XI102.XI1.MM1 N_XI0.XI102.NET6_XI0.XI102.XI1.MM1_d
+ N_MIN3_XI0.XI102.XI1.MM1_g N_VDD_XI0.XI102.XI1.MM1_s N_VDD_XI0.XI102.XI1.MM3_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.65e-13 PD=7.4e-07 PS=2.52e-06
mXI0.XI88.XI1.MM1 N_XI0.XI88.NET6_XI0.XI88.XI1.MM1_d N_MIN2_XI0.XI88.XI1.MM1_g
+ N_VDD_XI0.XI88.XI1.MM1_s N_VDD_XI0.XI88.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=5.55e-13 AS=7.65e-13 PD=7.4e-07 PS=2.52e-06
mXI0.XI82.XI1.MM1 N_XI0.XI82.NET6_XI0.XI82.XI1.MM1_d N_MIN1_XI0.XI82.XI1.MM1_g
+ N_VDD_XI0.XI82.XI1.MM1_s N_VDD_XI0.XI82.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=5.55e-13 AS=7.65e-13 PD=7.4e-07 PS=2.52e-06
mXI0.XI10.XI1.MM1 N_XI0.XI10.NET6_XI0.XI10.XI1.MM1_d N_MIN0_XI0.XI10.XI1.MM1_g
+ N_VDD_XI0.XI10.XI1.MM1_s N_VDD_XI0.XI10.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=5.55e-13 AS=7.65e-13 PD=7.4e-07 PS=2.52e-06
mXI0.XI134.MM5 N_XI0.XI134.NET25_XI0.XI134.MM5_d
+ N_XI0.XI134.NET43_XI0.XI134.MM5_g N_VDD_XI0.XI134.MM5_s
+ N_VDD_XI0.XI134.XI9.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=6.7125e-13 AS=9.675e-13
+ PD=8.95e-07 PS=2.79e-06
mXI0.XI153.XI0.MM1 N_XI0.G15_XI0.XI153.XI0.MM1_d
+ N_XI0.XI153.NET6_XI0.XI153.XI0.MM1_g N_VDD_XI0.XI153.XI0.MM1_s
+ N_VDD_XI0.XI153.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI0.XI154.XI0.MM1 N_XI0.G14_XI0.XI154.XI0.MM1_d
+ N_XI0.XI154.NET6_XI0.XI154.XI0.MM1_g N_VDD_XI0.XI154.XI0.MM1_s
+ N_VDD_XI0.XI154.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI0.XI157.XI0.MM1 N_XI0.G13_XI0.XI157.XI0.MM1_d
+ N_XI0.XI157.NET6_XI0.XI157.XI0.MM1_g N_VDD_XI0.XI157.XI0.MM1_s
+ N_VDD_XI0.XI157.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI0.XI156.XI0.MM1 N_XI0.G12_XI0.XI156.XI0.MM1_d
+ N_XI0.XI156.NET6_XI0.XI156.XI0.MM1_g N_VDD_XI0.XI156.XI0.MM1_s
+ N_VDD_XI0.XI156.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI0.XI155.XI0.MM1 N_XI0.G11_XI0.XI155.XI0.MM1_d
+ N_XI0.XI155.NET6_XI0.XI155.XI0.MM1_g N_VDD_XI0.XI155.XI0.MM1_s
+ N_VDD_XI0.XI155.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI0.XI133.XI0.MM1 N_XI0.G10_XI0.XI133.XI0.MM1_d
+ N_XI0.XI133.NET6_XI0.XI133.XI0.MM1_g N_VDD_XI0.XI133.XI0.MM1_s
+ N_VDD_XI0.XI133.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI0.XI132.XI0.MM1 N_XI0.G9_XI0.XI132.XI0.MM1_d
+ N_XI0.XI132.NET6_XI0.XI132.XI0.MM1_g N_VDD_XI0.XI132.XI0.MM1_s
+ N_VDD_XI0.XI132.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI0.XI131.XI0.MM1 N_XI0.G8_XI0.XI131.XI0.MM1_d
+ N_XI0.XI131.NET6_XI0.XI131.XI0.MM1_g N_VDD_XI0.XI131.XI0.MM1_s
+ N_VDD_XI0.XI131.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI0.XI111.XI0.MM1 N_XI0.G7_XI0.XI111.XI0.MM1_d
+ N_XI0.XI111.NET6_XI0.XI111.XI0.MM1_g N_VDD_XI0.XI111.XI0.MM1_s
+ N_VDD_XI0.XI111.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI0.XI110.XI0.MM1 N_XI0.G6_XI0.XI110.XI0.MM1_d
+ N_XI0.XI110.NET6_XI0.XI110.XI0.MM1_g N_VDD_XI0.XI110.XI0.MM1_s
+ N_VDD_XI0.XI110.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI0.XI103.XI0.MM1 N_XI0.G5_XI0.XI103.XI0.MM1_d
+ N_XI0.XI103.NET6_XI0.XI103.XI0.MM1_g N_VDD_XI0.XI103.XI0.MM1_s
+ N_VDD_XI0.XI103.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI0.XI102.XI0.MM1 N_XI0.G4_XI0.XI102.XI0.MM1_d
+ N_XI0.XI102.NET6_XI0.XI102.XI0.MM1_g N_VDD_XI0.XI102.XI0.MM1_s
+ N_VDD_XI0.XI102.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI0.XI88.XI0.MM1 N_XI0.G3_XI0.XI88.XI0.MM1_d N_XI0.XI88.NET6_XI0.XI88.XI0.MM1_g
+ N_VDD_XI0.XI88.XI0.MM1_s N_VDD_XI0.XI88.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI0.XI82.XI0.MM1 N_XI0.G2_XI0.XI82.XI0.MM1_d N_XI0.XI82.NET6_XI0.XI82.XI0.MM1_g
+ N_VDD_XI0.XI82.XI0.MM1_s N_VDD_XI0.XI82.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI0.XI10.XI0.MM1 N_XI0.G1_XI0.XI10.XI0.MM1_d N_XI0.XI10.NET6_XI0.XI10.XI0.MM1_g
+ N_VDD_XI0.XI10.XI0.MM1_s N_VDD_XI0.XI10.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI0.XI134.MM4 N_XI0.P16_XI0.XI134.MM4_d N_MIN15_XI0.XI134.MM4_g
+ N_XI0.XI134.NET25_XI0.XI134.MM4_s N_VDD_XI0.XI134.XI9.MM1_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.425e-12 AS=6.7125e-13 PD=1.9e-06 PS=8.95e-07
mXI0.XI137.XI9.MM1 N_XI0.XI137.NET43_XI0.XI137.XI9.MM1_d
+ N_NET595_XI0.XI137.XI9.MM1_g N_VDD_XI0.XI137.XI9.MM1_s
+ N_VDD_XI0.XI153.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI0.XI140.XI9.MM1 N_XI0.XI140.NET43_XI0.XI140.XI9.MM1_d
+ N_NET596_XI0.XI140.XI9.MM1_g N_VDD_XI0.XI140.XI9.MM1_s
+ N_VDD_XI0.XI154.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI0.XI149.XI9.MM1 N_XI0.XI149.NET43_XI0.XI149.XI9.MM1_d
+ N_NET597_XI0.XI149.XI9.MM1_g N_VDD_XI0.XI149.XI9.MM1_s
+ N_VDD_XI0.XI157.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI0.XI146.XI9.MM1 N_XI0.XI146.NET43_XI0.XI146.XI9.MM1_d
+ N_NET598_XI0.XI146.XI9.MM1_g N_VDD_XI0.XI146.XI9.MM1_s
+ N_VDD_XI0.XI156.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI0.XI143.XI9.MM1 N_XI0.XI143.NET43_XI0.XI143.XI9.MM1_d
+ N_NET599_XI0.XI143.XI9.MM1_g N_VDD_XI0.XI143.XI9.MM1_s
+ N_VDD_XI0.XI155.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI0.XI128.XI9.MM1 N_XI0.XI128.NET43_XI0.XI128.XI9.MM1_d
+ N_NET600_XI0.XI128.XI9.MM1_g N_VDD_XI0.XI128.XI9.MM1_s
+ N_VDD_XI0.XI133.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI0.XI125.XI9.MM1 N_XI0.XI125.NET43_XI0.XI125.XI9.MM1_d
+ N_NET601_XI0.XI125.XI9.MM1_g N_VDD_XI0.XI125.XI9.MM1_s
+ N_VDD_XI0.XI132.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI0.XI122.XI9.MM1 N_XI0.XI122.NET43_XI0.XI122.XI9.MM1_d
+ N_NET602_XI0.XI122.XI9.MM1_g N_VDD_XI0.XI122.XI9.MM1_s
+ N_VDD_XI0.XI131.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI0.XI114.XI9.MM1 N_XI0.XI114.NET43_XI0.XI114.XI9.MM1_d
+ N_NET603_XI0.XI114.XI9.MM1_g N_VDD_XI0.XI114.XI9.MM1_s
+ N_VDD_XI0.XI111.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI0.XI109.XI9.MM1 N_XI0.XI109.NET43_XI0.XI109.XI9.MM1_d
+ N_NET604_XI0.XI109.XI9.MM1_g N_VDD_XI0.XI109.XI9.MM1_s
+ N_VDD_XI0.XI110.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI0.XI106.XI9.MM1 N_XI0.XI106.NET43_XI0.XI106.XI9.MM1_d
+ N_NET605_XI0.XI106.XI9.MM1_g N_VDD_XI0.XI106.XI9.MM1_s
+ N_VDD_XI0.XI103.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI0.XI101.XI9.MM1 N_XI0.XI101.NET43_XI0.XI101.XI9.MM1_d
+ N_NET606_XI0.XI101.XI9.MM1_g N_VDD_XI0.XI101.XI9.MM1_s
+ N_VDD_XI0.XI102.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI0.XI86.XI9.MM1 N_XI0.XI86.NET43_XI0.XI86.XI9.MM1_d
+ N_NET607_XI0.XI86.XI9.MM1_g N_VDD_XI0.XI86.XI9.MM1_s N_VDD_XI0.XI88.XI1.MM3_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI0.XI80.XI9.MM1 N_XI0.XI80.NET43_XI0.XI80.XI9.MM1_d
+ N_NET608_XI0.XI80.XI9.MM1_g N_VDD_XI0.XI80.XI9.MM1_s N_VDD_XI0.XI82.XI1.MM3_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI0.XI26.XI9.MM1 N_XI0.XI26.NET43_XI0.XI26.XI9.MM1_d
+ N_NET609_XI0.XI26.XI9.MM1_g N_VDD_XI0.XI26.XI9.MM1_s N_VDD_XI0.XI10.XI1.MM3_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI0.XI134.MM3 N_XI0.P16_XI0.XI134.MM3_d N_XI0.XI134.NET39_XI0.XI134.MM3_g
+ N_XI0.XI134.NET37_XI0.XI134.MM3_s N_VDD_XI0.XI134.XI9.MM1_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.425e-12 AS=5.4375e-13 PD=1.9e-06 PS=7.25e-07
mXI0.XI134.MM1 N_XI0.XI134.NET37_XI0.XI134.MM1_d N_NET594_XI0.XI134.MM1_g
+ N_VDD_XI0.XI134.MM1_s N_VDD_XI0.XI134.XI9.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=5.4375e-13 AS=7.65e-13 PD=7.25e-07 PS=2.52e-06
mXI0.XI137.MM5 N_XI0.XI137.NET25_XI0.XI137.MM5_d
+ N_XI0.XI137.NET43_XI0.XI137.MM5_g N_VDD_XI0.XI137.MM5_s
+ N_VDD_XI0.XI153.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=6.7125e-13 AS=9.675e-13
+ PD=8.95e-07 PS=2.79e-06
mXI0.XI140.MM5 N_XI0.XI140.NET25_XI0.XI140.MM5_d
+ N_XI0.XI140.NET43_XI0.XI140.MM5_g N_VDD_XI0.XI140.MM5_s
+ N_VDD_XI0.XI154.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=6.7125e-13 AS=9.675e-13
+ PD=8.95e-07 PS=2.79e-06
mXI0.XI149.MM5 N_XI0.XI149.NET25_XI0.XI149.MM5_d
+ N_XI0.XI149.NET43_XI0.XI149.MM5_g N_VDD_XI0.XI149.MM5_s
+ N_VDD_XI0.XI157.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=6.7125e-13 AS=9.675e-13
+ PD=8.95e-07 PS=2.79e-06
mXI0.XI146.MM5 N_XI0.XI146.NET25_XI0.XI146.MM5_d
+ N_XI0.XI146.NET43_XI0.XI146.MM5_g N_VDD_XI0.XI146.MM5_s
+ N_VDD_XI0.XI156.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=6.7125e-13 AS=9.675e-13
+ PD=8.95e-07 PS=2.79e-06
mXI0.XI143.MM5 N_XI0.XI143.NET25_XI0.XI143.MM5_d
+ N_XI0.XI143.NET43_XI0.XI143.MM5_g N_VDD_XI0.XI143.MM5_s
+ N_VDD_XI0.XI155.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=6.7125e-13 AS=9.675e-13
+ PD=8.95e-07 PS=2.79e-06
mXI0.XI128.MM5 N_XI0.XI128.NET25_XI0.XI128.MM5_d
+ N_XI0.XI128.NET43_XI0.XI128.MM5_g N_VDD_XI0.XI128.MM5_s
+ N_VDD_XI0.XI133.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=6.7125e-13 AS=9.675e-13
+ PD=8.95e-07 PS=2.79e-06
mXI0.XI125.MM5 N_XI0.XI125.NET25_XI0.XI125.MM5_d
+ N_XI0.XI125.NET43_XI0.XI125.MM5_g N_VDD_XI0.XI125.MM5_s
+ N_VDD_XI0.XI132.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=6.7125e-13 AS=9.675e-13
+ PD=8.95e-07 PS=2.79e-06
mXI0.XI122.MM5 N_XI0.XI122.NET25_XI0.XI122.MM5_d
+ N_XI0.XI122.NET43_XI0.XI122.MM5_g N_VDD_XI0.XI122.MM5_s
+ N_VDD_XI0.XI131.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=6.7125e-13 AS=9.675e-13
+ PD=8.95e-07 PS=2.79e-06
mXI0.XI114.MM5 N_XI0.XI114.NET25_XI0.XI114.MM5_d
+ N_XI0.XI114.NET43_XI0.XI114.MM5_g N_VDD_XI0.XI114.MM5_s
+ N_VDD_XI0.XI111.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=6.7125e-13 AS=9.675e-13
+ PD=8.95e-07 PS=2.79e-06
mXI0.XI109.MM5 N_XI0.XI109.NET25_XI0.XI109.MM5_d
+ N_XI0.XI109.NET43_XI0.XI109.MM5_g N_VDD_XI0.XI109.MM5_s
+ N_VDD_XI0.XI110.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=6.7125e-13 AS=9.675e-13
+ PD=8.95e-07 PS=2.79e-06
mXI0.XI106.MM5 N_XI0.XI106.NET25_XI0.XI106.MM5_d
+ N_XI0.XI106.NET43_XI0.XI106.MM5_g N_VDD_XI0.XI106.MM5_s
+ N_VDD_XI0.XI103.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=6.7125e-13 AS=9.675e-13
+ PD=8.95e-07 PS=2.79e-06
mXI0.XI101.MM5 N_XI0.XI101.NET25_XI0.XI101.MM5_d
+ N_XI0.XI101.NET43_XI0.XI101.MM5_g N_VDD_XI0.XI101.MM5_s
+ N_VDD_XI0.XI102.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=6.7125e-13 AS=9.675e-13
+ PD=8.95e-07 PS=2.79e-06
mXI0.XI86.MM5 N_XI0.XI86.NET25_XI0.XI86.MM5_d N_XI0.XI86.NET43_XI0.XI86.MM5_g
+ N_VDD_XI0.XI86.MM5_s N_VDD_XI0.XI88.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=6.7125e-13 AS=9.675e-13 PD=8.95e-07 PS=2.79e-06
mXI0.XI80.MM5 N_XI0.XI80.NET25_XI0.XI80.MM5_d N_XI0.XI80.NET43_XI0.XI80.MM5_g
+ N_VDD_XI0.XI80.MM5_s N_VDD_XI0.XI82.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=6.7125e-13 AS=9.675e-13 PD=8.95e-07 PS=2.79e-06
mXI0.XI26.MM5 N_XI0.XI26.NET25_XI0.XI26.MM5_d N_XI0.XI26.NET43_XI0.XI26.MM5_g
+ N_VDD_XI0.XI26.MM5_s N_VDD_XI0.XI10.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=6.7125e-13 AS=9.675e-13 PD=8.95e-07 PS=2.79e-06
mXI0.XI137.MM4 N_XI0.P15_XI0.XI137.MM4_d N_MIN14_XI0.XI137.MM4_g
+ N_XI0.XI137.NET25_XI0.XI137.MM4_s N_VDD_XI0.XI153.XI1.MM3_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.425e-12 AS=6.7125e-13 PD=1.9e-06 PS=8.95e-07
mXI0.XI140.MM4 N_XI0.P14_XI0.XI140.MM4_d N_MIN13_XI0.XI140.MM4_g
+ N_XI0.XI140.NET25_XI0.XI140.MM4_s N_VDD_XI0.XI154.XI1.MM3_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.425e-12 AS=6.7125e-13 PD=1.9e-06 PS=8.95e-07
mXI0.XI149.MM4 N_XI0.P13_XI0.XI149.MM4_d N_MIN12_XI0.XI149.MM4_g
+ N_XI0.XI149.NET25_XI0.XI149.MM4_s N_VDD_XI0.XI157.XI1.MM3_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.425e-12 AS=6.7125e-13 PD=1.9e-06 PS=8.95e-07
mXI0.XI146.MM4 N_XI0.P12_XI0.XI146.MM4_d N_MIN11_XI0.XI146.MM4_g
+ N_XI0.XI146.NET25_XI0.XI146.MM4_s N_VDD_XI0.XI156.XI1.MM3_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.425e-12 AS=6.7125e-13 PD=1.9e-06 PS=8.95e-07
mXI0.XI143.MM4 N_XI0.P11_XI0.XI143.MM4_d N_MIN10_XI0.XI143.MM4_g
+ N_XI0.XI143.NET25_XI0.XI143.MM4_s N_VDD_XI0.XI155.XI1.MM3_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.425e-12 AS=6.7125e-13 PD=1.9e-06 PS=8.95e-07
mXI0.XI128.MM4 N_XI0.P10_XI0.XI128.MM4_d N_MIN9_XI0.XI128.MM4_g
+ N_XI0.XI128.NET25_XI0.XI128.MM4_s N_VDD_XI0.XI133.XI1.MM3_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.425e-12 AS=6.7125e-13 PD=1.9e-06 PS=8.95e-07
mXI0.XI125.MM4 N_XI0.P9_XI0.XI125.MM4_d N_MIN8_XI0.XI125.MM4_g
+ N_XI0.XI125.NET25_XI0.XI125.MM4_s N_VDD_XI0.XI132.XI1.MM3_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.425e-12 AS=6.7125e-13 PD=1.9e-06 PS=8.95e-07
mXI0.XI122.MM4 N_XI0.P8_XI0.XI122.MM4_d N_MIN7_XI0.XI122.MM4_g
+ N_XI0.XI122.NET25_XI0.XI122.MM4_s N_VDD_XI0.XI131.XI1.MM3_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.425e-12 AS=6.7125e-13 PD=1.9e-06 PS=8.95e-07
mXI0.XI114.MM4 N_XI0.P7_XI0.XI114.MM4_d N_MIN6_XI0.XI114.MM4_g
+ N_XI0.XI114.NET25_XI0.XI114.MM4_s N_VDD_XI0.XI111.XI1.MM3_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.425e-12 AS=6.7125e-13 PD=1.9e-06 PS=8.95e-07
mXI0.XI109.MM4 N_XI0.P6_XI0.XI109.MM4_d N_MIN5_XI0.XI109.MM4_g
+ N_XI0.XI109.NET25_XI0.XI109.MM4_s N_VDD_XI0.XI110.XI1.MM3_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.425e-12 AS=6.7125e-13 PD=1.9e-06 PS=8.95e-07
mXI0.XI106.MM4 N_XI0.P5_XI0.XI106.MM4_d N_MIN4_XI0.XI106.MM4_g
+ N_XI0.XI106.NET25_XI0.XI106.MM4_s N_VDD_XI0.XI103.XI1.MM3_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.425e-12 AS=6.7125e-13 PD=1.9e-06 PS=8.95e-07
mXI0.XI101.MM4 N_XI0.P4_XI0.XI101.MM4_d N_MIN3_XI0.XI101.MM4_g
+ N_XI0.XI101.NET25_XI0.XI101.MM4_s N_VDD_XI0.XI102.XI1.MM3_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.425e-12 AS=6.7125e-13 PD=1.9e-06 PS=8.95e-07
mXI0.XI86.MM4 N_XI0.P3_XI0.XI86.MM4_d N_MIN2_XI0.XI86.MM4_g
+ N_XI0.XI86.NET25_XI0.XI86.MM4_s N_VDD_XI0.XI88.XI1.MM3_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.425e-12 AS=6.7125e-13 PD=1.9e-06 PS=8.95e-07
mXI0.XI80.MM4 N_XI0.P2_XI0.XI80.MM4_d N_MIN1_XI0.XI80.MM4_g
+ N_XI0.XI80.NET25_XI0.XI80.MM4_s N_VDD_XI0.XI82.XI1.MM3_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.425e-12 AS=6.7125e-13 PD=1.9e-06 PS=8.95e-07
mXI0.XI26.MM4 N_XI0.P1_XI0.XI26.MM4_d N_MIN0_XI0.XI26.MM4_g
+ N_XI0.XI26.NET25_XI0.XI26.MM4_s N_VDD_XI0.XI10.XI1.MM3_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.425e-12 AS=6.7125e-13 PD=1.9e-06 PS=8.95e-07
mXI0.XI134.XI4.MM1 N_XI0.XI134.NET39_XI0.XI134.XI4.MM1_d
+ N_MIN15_XI0.XI134.XI4.MM1_g N_VDD_XI0.XI134.XI4.MM1_s
+ N_VDD_XI0.XI134.XI9.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI0.XI137.MM3 N_XI0.P15_XI0.XI137.MM3_d N_XI0.XI137.NET39_XI0.XI137.MM3_g
+ N_XI0.XI137.NET37_XI0.XI137.MM3_s N_VDD_XI0.XI153.XI1.MM3_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.425e-12 AS=5.4375e-13 PD=1.9e-06 PS=7.25e-07
mXI0.XI140.MM3 N_XI0.P14_XI0.XI140.MM3_d N_XI0.XI140.NET39_XI0.XI140.MM3_g
+ N_XI0.XI140.NET37_XI0.XI140.MM3_s N_VDD_XI0.XI154.XI1.MM3_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.425e-12 AS=5.4375e-13 PD=1.9e-06 PS=7.25e-07
mXI0.XI149.MM3 N_XI0.P13_XI0.XI149.MM3_d N_XI0.XI149.NET39_XI0.XI149.MM3_g
+ N_XI0.XI149.NET37_XI0.XI149.MM3_s N_VDD_XI0.XI157.XI1.MM3_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.425e-12 AS=5.4375e-13 PD=1.9e-06 PS=7.25e-07
mXI0.XI146.MM3 N_XI0.P12_XI0.XI146.MM3_d N_XI0.XI146.NET39_XI0.XI146.MM3_g
+ N_XI0.XI146.NET37_XI0.XI146.MM3_s N_VDD_XI0.XI156.XI1.MM3_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.425e-12 AS=5.4375e-13 PD=1.9e-06 PS=7.25e-07
mXI0.XI143.MM3 N_XI0.P11_XI0.XI143.MM3_d N_XI0.XI143.NET39_XI0.XI143.MM3_g
+ N_XI0.XI143.NET37_XI0.XI143.MM3_s N_VDD_XI0.XI155.XI1.MM3_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.425e-12 AS=5.4375e-13 PD=1.9e-06 PS=7.25e-07
mXI0.XI128.MM3 N_XI0.P10_XI0.XI128.MM3_d N_XI0.XI128.NET39_XI0.XI128.MM3_g
+ N_XI0.XI128.NET37_XI0.XI128.MM3_s N_VDD_XI0.XI133.XI1.MM3_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.425e-12 AS=5.4375e-13 PD=1.9e-06 PS=7.25e-07
mXI0.XI125.MM3 N_XI0.P9_XI0.XI125.MM3_d N_XI0.XI125.NET39_XI0.XI125.MM3_g
+ N_XI0.XI125.NET37_XI0.XI125.MM3_s N_VDD_XI0.XI132.XI1.MM3_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.425e-12 AS=5.4375e-13 PD=1.9e-06 PS=7.25e-07
mXI0.XI122.MM3 N_XI0.P8_XI0.XI122.MM3_d N_XI0.XI122.NET39_XI0.XI122.MM3_g
+ N_XI0.XI122.NET37_XI0.XI122.MM3_s N_VDD_XI0.XI131.XI1.MM3_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.425e-12 AS=5.4375e-13 PD=1.9e-06 PS=7.25e-07
mXI0.XI114.MM3 N_XI0.P7_XI0.XI114.MM3_d N_XI0.XI114.NET39_XI0.XI114.MM3_g
+ N_XI0.XI114.NET37_XI0.XI114.MM3_s N_VDD_XI0.XI111.XI1.MM3_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.425e-12 AS=5.4375e-13 PD=1.9e-06 PS=7.25e-07
mXI0.XI109.MM3 N_XI0.P6_XI0.XI109.MM3_d N_XI0.XI109.NET39_XI0.XI109.MM3_g
+ N_XI0.XI109.NET37_XI0.XI109.MM3_s N_VDD_XI0.XI110.XI1.MM3_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.425e-12 AS=5.4375e-13 PD=1.9e-06 PS=7.25e-07
mXI0.XI106.MM3 N_XI0.P5_XI0.XI106.MM3_d N_XI0.XI106.NET39_XI0.XI106.MM3_g
+ N_XI0.XI106.NET37_XI0.XI106.MM3_s N_VDD_XI0.XI103.XI1.MM3_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.425e-12 AS=5.4375e-13 PD=1.9e-06 PS=7.25e-07
mXI0.XI101.MM3 N_XI0.P4_XI0.XI101.MM3_d N_XI0.XI101.NET39_XI0.XI101.MM3_g
+ N_XI0.XI101.NET37_XI0.XI101.MM3_s N_VDD_XI0.XI102.XI1.MM3_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.425e-12 AS=5.4375e-13 PD=1.9e-06 PS=7.25e-07
mXI0.XI86.MM3 N_XI0.P3_XI0.XI86.MM3_d N_XI0.XI86.NET39_XI0.XI86.MM3_g
+ N_XI0.XI86.NET37_XI0.XI86.MM3_s N_VDD_XI0.XI88.XI1.MM3_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.425e-12 AS=5.4375e-13 PD=1.9e-06 PS=7.25e-07
mXI0.XI80.MM3 N_XI0.P2_XI0.XI80.MM3_d N_XI0.XI80.NET39_XI0.XI80.MM3_g
+ N_XI0.XI80.NET37_XI0.XI80.MM3_s N_VDD_XI0.XI82.XI1.MM3_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.425e-12 AS=5.4375e-13 PD=1.9e-06 PS=7.25e-07
mXI0.XI26.MM3 N_XI0.P1_XI0.XI26.MM3_d N_XI0.XI26.NET39_XI0.XI26.MM3_g
+ N_XI0.XI26.NET37_XI0.XI26.MM3_s N_VDD_XI0.XI10.XI1.MM3_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.425e-12 AS=5.4375e-13 PD=1.9e-06 PS=7.25e-07
mXI0.XI137.MM1 N_XI0.XI137.NET37_XI0.XI137.MM1_d N_NET595_XI0.XI137.MM1_g
+ N_VDD_XI0.XI137.MM1_s N_VDD_XI0.XI153.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=5.4375e-13 AS=7.65e-13 PD=7.25e-07 PS=2.52e-06
mXI0.XI140.MM1 N_XI0.XI140.NET37_XI0.XI140.MM1_d N_NET596_XI0.XI140.MM1_g
+ N_VDD_XI0.XI140.MM1_s N_VDD_XI0.XI154.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=5.4375e-13 AS=7.65e-13 PD=7.25e-07 PS=2.52e-06
mXI0.XI149.MM1 N_XI0.XI149.NET37_XI0.XI149.MM1_d N_NET597_XI0.XI149.MM1_g
+ N_VDD_XI0.XI149.MM1_s N_VDD_XI0.XI157.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=5.4375e-13 AS=7.65e-13 PD=7.25e-07 PS=2.52e-06
mXI0.XI146.MM1 N_XI0.XI146.NET37_XI0.XI146.MM1_d N_NET598_XI0.XI146.MM1_g
+ N_VDD_XI0.XI146.MM1_s N_VDD_XI0.XI156.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=5.4375e-13 AS=7.65e-13 PD=7.25e-07 PS=2.52e-06
mXI0.XI143.MM1 N_XI0.XI143.NET37_XI0.XI143.MM1_d N_NET599_XI0.XI143.MM1_g
+ N_VDD_XI0.XI143.MM1_s N_VDD_XI0.XI155.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=5.4375e-13 AS=7.65e-13 PD=7.25e-07 PS=2.52e-06
mXI0.XI128.MM1 N_XI0.XI128.NET37_XI0.XI128.MM1_d N_NET600_XI0.XI128.MM1_g
+ N_VDD_XI0.XI128.MM1_s N_VDD_XI0.XI133.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=5.4375e-13 AS=7.65e-13 PD=7.25e-07 PS=2.52e-06
mXI0.XI125.MM1 N_XI0.XI125.NET37_XI0.XI125.MM1_d N_NET601_XI0.XI125.MM1_g
+ N_VDD_XI0.XI125.MM1_s N_VDD_XI0.XI132.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=5.4375e-13 AS=7.65e-13 PD=7.25e-07 PS=2.52e-06
mXI0.XI122.MM1 N_XI0.XI122.NET37_XI0.XI122.MM1_d N_NET602_XI0.XI122.MM1_g
+ N_VDD_XI0.XI122.MM1_s N_VDD_XI0.XI131.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=5.4375e-13 AS=7.65e-13 PD=7.25e-07 PS=2.52e-06
mXI0.XI114.MM1 N_XI0.XI114.NET37_XI0.XI114.MM1_d N_NET603_XI0.XI114.MM1_g
+ N_VDD_XI0.XI114.MM1_s N_VDD_XI0.XI111.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=5.4375e-13 AS=7.65e-13 PD=7.25e-07 PS=2.52e-06
mXI0.XI109.MM1 N_XI0.XI109.NET37_XI0.XI109.MM1_d N_NET604_XI0.XI109.MM1_g
+ N_VDD_XI0.XI109.MM1_s N_VDD_XI0.XI110.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=5.4375e-13 AS=7.65e-13 PD=7.25e-07 PS=2.52e-06
mXI0.XI106.MM1 N_XI0.XI106.NET37_XI0.XI106.MM1_d N_NET605_XI0.XI106.MM1_g
+ N_VDD_XI0.XI106.MM1_s N_VDD_XI0.XI103.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=5.4375e-13 AS=7.65e-13 PD=7.25e-07 PS=2.52e-06
mXI0.XI101.MM1 N_XI0.XI101.NET37_XI0.XI101.MM1_d N_NET606_XI0.XI101.MM1_g
+ N_VDD_XI0.XI101.MM1_s N_VDD_XI0.XI102.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=5.4375e-13 AS=7.65e-13 PD=7.25e-07 PS=2.52e-06
mXI0.XI86.MM1 N_XI0.XI86.NET37_XI0.XI86.MM1_d N_NET607_XI0.XI86.MM1_g
+ N_VDD_XI0.XI86.MM1_s N_VDD_XI0.XI88.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=5.4375e-13 AS=7.65e-13 PD=7.25e-07 PS=2.52e-06
mXI0.XI80.MM1 N_XI0.XI80.NET37_XI0.XI80.MM1_d N_NET608_XI0.XI80.MM1_g
+ N_VDD_XI0.XI80.MM1_s N_VDD_XI0.XI82.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=5.4375e-13 AS=7.65e-13 PD=7.25e-07 PS=2.52e-06
mXI0.XI26.MM1 N_XI0.XI26.NET37_XI0.XI26.MM1_d N_NET609_XI0.XI26.MM1_g
+ N_VDD_XI0.XI26.MM1_s N_VDD_XI0.XI10.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=5.4375e-13 AS=7.65e-13 PD=7.25e-07 PS=2.52e-06
mXI0.XI182.XI9.MM1 N_XI0.XI182.NET43_XI0.XI182.XI9.MM1_d
+ N_XI0.P16_XI0.XI182.XI9.MM1_g N_VDD_XI0.XI182.XI9.MM1_s
+ N_VDD_XI0.XI134.XI9.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI0.XI137.XI4.MM1 N_XI0.XI137.NET39_XI0.XI137.XI4.MM1_d
+ N_MIN14_XI0.XI137.XI4.MM1_g N_VDD_XI0.XI137.XI4.MM1_s
+ N_VDD_XI0.XI153.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI0.XI140.XI4.MM1 N_XI0.XI140.NET39_XI0.XI140.XI4.MM1_d
+ N_MIN13_XI0.XI140.XI4.MM1_g N_VDD_XI0.XI140.XI4.MM1_s
+ N_VDD_XI0.XI154.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI0.XI149.XI4.MM1 N_XI0.XI149.NET39_XI0.XI149.XI4.MM1_d
+ N_MIN12_XI0.XI149.XI4.MM1_g N_VDD_XI0.XI149.XI4.MM1_s
+ N_VDD_XI0.XI157.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI0.XI146.XI4.MM1 N_XI0.XI146.NET39_XI0.XI146.XI4.MM1_d
+ N_MIN11_XI0.XI146.XI4.MM1_g N_VDD_XI0.XI146.XI4.MM1_s
+ N_VDD_XI0.XI156.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI0.XI143.XI4.MM1 N_XI0.XI143.NET39_XI0.XI143.XI4.MM1_d
+ N_MIN10_XI0.XI143.XI4.MM1_g N_VDD_XI0.XI143.XI4.MM1_s
+ N_VDD_XI0.XI155.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI0.XI128.XI4.MM1 N_XI0.XI128.NET39_XI0.XI128.XI4.MM1_d
+ N_MIN9_XI0.XI128.XI4.MM1_g N_VDD_XI0.XI128.XI4.MM1_s N_VDD_XI0.XI133.XI1.MM3_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI0.XI125.XI4.MM1 N_XI0.XI125.NET39_XI0.XI125.XI4.MM1_d
+ N_MIN8_XI0.XI125.XI4.MM1_g N_VDD_XI0.XI125.XI4.MM1_s N_VDD_XI0.XI132.XI1.MM3_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI0.XI122.XI4.MM1 N_XI0.XI122.NET39_XI0.XI122.XI4.MM1_d
+ N_MIN7_XI0.XI122.XI4.MM1_g N_VDD_XI0.XI122.XI4.MM1_s N_VDD_XI0.XI131.XI1.MM3_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI0.XI114.XI4.MM1 N_XI0.XI114.NET39_XI0.XI114.XI4.MM1_d
+ N_MIN6_XI0.XI114.XI4.MM1_g N_VDD_XI0.XI114.XI4.MM1_s N_VDD_XI0.XI111.XI1.MM3_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI0.XI109.XI4.MM1 N_XI0.XI109.NET39_XI0.XI109.XI4.MM1_d
+ N_MIN5_XI0.XI109.XI4.MM1_g N_VDD_XI0.XI109.XI4.MM1_s N_VDD_XI0.XI110.XI1.MM3_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI0.XI106.XI4.MM1 N_XI0.XI106.NET39_XI0.XI106.XI4.MM1_d
+ N_MIN4_XI0.XI106.XI4.MM1_g N_VDD_XI0.XI106.XI4.MM1_s N_VDD_XI0.XI103.XI1.MM3_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI0.XI101.XI4.MM1 N_XI0.XI101.NET39_XI0.XI101.XI4.MM1_d
+ N_MIN3_XI0.XI101.XI4.MM1_g N_VDD_XI0.XI101.XI4.MM1_s N_VDD_XI0.XI102.XI1.MM3_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI0.XI86.XI4.MM1 N_XI0.XI86.NET39_XI0.XI86.XI4.MM1_d N_MIN2_XI0.XI86.XI4.MM1_g
+ N_VDD_XI0.XI86.XI4.MM1_s N_VDD_XI0.XI88.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI0.XI80.XI4.MM1 N_XI0.XI80.NET39_XI0.XI80.XI4.MM1_d N_MIN1_XI0.XI80.XI4.MM1_g
+ N_VDD_XI0.XI80.XI4.MM1_s N_VDD_XI0.XI82.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI0.XI26.XI4.MM1 N_XI0.XI26.NET39_XI0.XI26.XI4.MM1_d N_MIN0_XI0.XI26.XI4.MM1_g
+ N_VDD_XI0.XI26.XI4.MM1_s N_VDD_XI0.XI10.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI0.XI182.MM5 N_XI0.XI182.NET25_XI0.XI182.MM5_d
+ N_XI0.XI182.NET43_XI0.XI182.MM5_g N_VDD_XI0.XI182.MM5_s
+ N_VDD_XI0.XI134.XI9.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=6.7125e-13 AS=9.675e-13
+ PD=8.95e-07 PS=2.79e-06
mXI0.XI168.XI1.XI1.MM1 N_XI0.XI168.XI1.NET6_XI0.XI168.XI1.XI1.MM1_d
+ N_XI0.NET288_XI0.XI168.XI1.XI1.MM1_g N_VDD_XI0.XI168.XI1.XI1.MM1_s
+ N_VDD_XI0.XI153.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.35e-13
+ PD=7.4e-07 PS=2.48e-06
mXI0.XI167.XI1.XI1.MM1 N_XI0.XI167.XI1.NET6_XI0.XI167.XI1.XI1.MM1_d
+ N_XI0.NET282_XI0.XI167.XI1.XI1.MM1_g N_VDD_XI0.XI167.XI1.XI1.MM1_s
+ N_VDD_XI0.XI154.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.35e-13
+ PD=7.4e-07 PS=2.48e-06
mXI0.XI166.XI1.XI1.MM1 N_XI0.XI166.XI1.NET6_XI0.XI166.XI1.XI1.MM1_d
+ N_XI0.NET276_XI0.XI166.XI1.XI1.MM1_g N_VDD_XI0.XI166.XI1.XI1.MM1_s
+ N_VDD_XI0.XI157.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.35e-13
+ PD=7.4e-07 PS=2.48e-06
mXI0.XI165.XI1.XI1.MM1 N_XI0.XI165.XI1.NET6_XI0.XI165.XI1.XI1.MM1_d
+ N_XI0.NET270_XI0.XI165.XI1.XI1.MM1_g N_VDD_XI0.XI165.XI1.XI1.MM1_s
+ N_VDD_XI0.XI156.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.35e-13
+ PD=7.4e-07 PS=2.48e-06
mXI0.XI159.XI1.XI1.MM1 N_XI0.XI159.XI1.NET6_XI0.XI159.XI1.XI1.MM1_d
+ N_XI0.NET246_XI0.XI159.XI1.XI1.MM1_g N_VDD_XI0.XI159.XI1.XI1.MM1_s
+ N_VDD_XI0.XI155.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.35e-13
+ PD=7.4e-07 PS=2.48e-06
mXI0.XI160.XI1.XI1.MM1 N_XI0.XI160.XI1.NET6_XI0.XI160.XI1.XI1.MM1_d
+ N_XI0.NET252_XI0.XI160.XI1.XI1.MM1_g N_VDD_XI0.XI160.XI1.XI1.MM1_s
+ N_VDD_XI0.XI133.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.35e-13
+ PD=7.4e-07 PS=2.48e-06
mXI0.XI161.XI1.XI1.MM1 N_XI0.XI161.XI1.NET6_XI0.XI161.XI1.XI1.MM1_d
+ N_XI0.NET258_XI0.XI161.XI1.XI1.MM1_g N_VDD_XI0.XI161.XI1.XI1.MM1_s
+ N_VDD_XI0.XI132.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.35e-13
+ PD=7.4e-07 PS=2.48e-06
mXI0.XI162.XI1.XI1.MM1 N_XI0.XI162.XI1.NET6_XI0.XI162.XI1.XI1.MM1_d
+ N_XI0.NET264_XI0.XI162.XI1.XI1.MM1_g N_VDD_XI0.XI162.XI1.XI1.MM1_s
+ N_VDD_XI0.XI131.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.35e-13
+ PD=7.4e-07 PS=2.48e-06
mXI0.XI121.XI1.XI1.MM1 N_XI0.XI121.XI1.NET6_XI0.XI121.XI1.XI1.MM1_d
+ N_XI0.NET204_XI0.XI121.XI1.XI1.MM1_g N_VDD_XI0.XI121.XI1.XI1.MM1_s
+ N_VDD_XI0.XI111.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.35e-13
+ PD=7.4e-07 PS=2.48e-06
mXI0.XI120.XI1.XI1.MM1 N_XI0.XI120.XI1.NET6_XI0.XI120.XI1.XI1.MM1_d
+ N_XI0.NET210_XI0.XI120.XI1.XI1.MM1_g N_VDD_XI0.XI120.XI1.XI1.MM1_s
+ N_VDD_XI0.XI110.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.35e-13
+ PD=7.4e-07 PS=2.48e-06
mXI0.XI119.XI1.XI1.MM1 N_XI0.XI119.XI1.NET6_XI0.XI119.XI1.XI1.MM1_d
+ N_XI0.NET216_XI0.XI119.XI1.XI1.MM1_g N_VDD_XI0.XI119.XI1.XI1.MM1_s
+ N_VDD_XI0.XI103.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.35e-13
+ PD=7.4e-07 PS=2.48e-06
mXI0.XI118.XI1.XI1.MM1 N_XI0.XI118.XI1.NET6_XI0.XI118.XI1.XI1.MM1_d
+ N_XI0.NET222_XI0.XI118.XI1.XI1.MM1_g N_VDD_XI0.XI118.XI1.XI1.MM1_s
+ N_VDD_XI0.XI102.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.35e-13
+ PD=7.4e-07 PS=2.48e-06
mXI0.XI91.XI1.XI1.MM1 N_XI0.XI91.XI1.NET6_XI0.XI91.XI1.XI1.MM1_d
+ N_XI0.NET228_XI0.XI91.XI1.XI1.MM1_g N_VDD_XI0.XI91.XI1.XI1.MM1_s
+ N_VDD_XI0.XI88.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.35e-13
+ PD=7.4e-07 PS=2.48e-06
mXI0.XI90.XI1.XI1.MM1 N_XI0.XI90.XI1.NET6_XI0.XI90.XI1.XI1.MM1_d
+ N_XI0.NET240_XI0.XI90.XI1.XI1.MM1_g N_VDD_XI0.XI90.XI1.XI1.MM1_s
+ N_VDD_XI0.XI82.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.35e-13
+ PD=7.4e-07 PS=2.48e-06
mXI0.XI89.XI1.XI1.MM1 N_XI0.XI89.XI1.NET6_XI0.XI89.XI1.XI1.MM1_d
+ N_CIN2_XI0.XI89.XI1.XI1.MM1_g N_VDD_XI0.XI89.XI1.XI1.MM1_s
+ N_VDD_XI0.XI10.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.35e-13
+ PD=7.4e-07 PS=2.48e-06
mXI0.XI182.MM4 N_NET141_XI0.XI182.MM4_d N_XI0.NET198_XI0.XI182.MM4_g
+ N_XI0.XI182.NET25_XI0.XI182.MM4_s N_VDD_XI0.XI134.XI9.MM1_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.425e-12 AS=6.7125e-13 PD=1.9e-06 PS=8.95e-07
mXI0.XI168.XI1.XI1.MM3 N_XI0.XI168.XI1.NET6_XI0.XI168.XI1.XI1.MM3_d
+ N_XI0.P15_XI0.XI168.XI1.XI1.MM3_g N_VDD_XI0.XI168.XI1.XI1.MM3_s
+ N_VDD_XI0.XI153.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.65e-13
+ PD=7.4e-07 PS=2.52e-06
mXI0.XI167.XI1.XI1.MM3 N_XI0.XI167.XI1.NET6_XI0.XI167.XI1.XI1.MM3_d
+ N_XI0.P14_XI0.XI167.XI1.XI1.MM3_g N_VDD_XI0.XI167.XI1.XI1.MM3_s
+ N_VDD_XI0.XI154.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.65e-13
+ PD=7.4e-07 PS=2.52e-06
mXI0.XI166.XI1.XI1.MM3 N_XI0.XI166.XI1.NET6_XI0.XI166.XI1.XI1.MM3_d
+ N_XI0.P13_XI0.XI166.XI1.XI1.MM3_g N_VDD_XI0.XI166.XI1.XI1.MM3_s
+ N_VDD_XI0.XI157.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.65e-13
+ PD=7.4e-07 PS=2.52e-06
mXI0.XI165.XI1.XI1.MM3 N_XI0.XI165.XI1.NET6_XI0.XI165.XI1.XI1.MM3_d
+ N_XI0.P12_XI0.XI165.XI1.XI1.MM3_g N_VDD_XI0.XI165.XI1.XI1.MM3_s
+ N_VDD_XI0.XI156.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.65e-13
+ PD=7.4e-07 PS=2.52e-06
mXI0.XI159.XI1.XI1.MM3 N_XI0.XI159.XI1.NET6_XI0.XI159.XI1.XI1.MM3_d
+ N_XI0.P11_XI0.XI159.XI1.XI1.MM3_g N_VDD_XI0.XI159.XI1.XI1.MM3_s
+ N_VDD_XI0.XI155.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.65e-13
+ PD=7.4e-07 PS=2.52e-06
mXI0.XI160.XI1.XI1.MM3 N_XI0.XI160.XI1.NET6_XI0.XI160.XI1.XI1.MM3_d
+ N_XI0.P10_XI0.XI160.XI1.XI1.MM3_g N_VDD_XI0.XI160.XI1.XI1.MM3_s
+ N_VDD_XI0.XI133.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.65e-13
+ PD=7.4e-07 PS=2.52e-06
mXI0.XI161.XI1.XI1.MM3 N_XI0.XI161.XI1.NET6_XI0.XI161.XI1.XI1.MM3_d
+ N_XI0.P9_XI0.XI161.XI1.XI1.MM3_g N_VDD_XI0.XI161.XI1.XI1.MM3_s
+ N_VDD_XI0.XI132.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.65e-13
+ PD=7.4e-07 PS=2.52e-06
mXI0.XI162.XI1.XI1.MM3 N_XI0.XI162.XI1.NET6_XI0.XI162.XI1.XI1.MM3_d
+ N_XI0.P8_XI0.XI162.XI1.XI1.MM3_g N_VDD_XI0.XI162.XI1.XI1.MM3_s
+ N_VDD_XI0.XI131.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.65e-13
+ PD=7.4e-07 PS=2.52e-06
mXI0.XI121.XI1.XI1.MM3 N_XI0.XI121.XI1.NET6_XI0.XI121.XI1.XI1.MM3_d
+ N_XI0.P7_XI0.XI121.XI1.XI1.MM3_g N_VDD_XI0.XI121.XI1.XI1.MM3_s
+ N_VDD_XI0.XI111.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.65e-13
+ PD=7.4e-07 PS=2.52e-06
mXI0.XI120.XI1.XI1.MM3 N_XI0.XI120.XI1.NET6_XI0.XI120.XI1.XI1.MM3_d
+ N_XI0.P6_XI0.XI120.XI1.XI1.MM3_g N_VDD_XI0.XI120.XI1.XI1.MM3_s
+ N_VDD_XI0.XI110.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.65e-13
+ PD=7.4e-07 PS=2.52e-06
mXI0.XI119.XI1.XI1.MM3 N_XI0.XI119.XI1.NET6_XI0.XI119.XI1.XI1.MM3_d
+ N_XI0.P5_XI0.XI119.XI1.XI1.MM3_g N_VDD_XI0.XI119.XI1.XI1.MM3_s
+ N_VDD_XI0.XI103.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.65e-13
+ PD=7.4e-07 PS=2.52e-06
mXI0.XI118.XI1.XI1.MM3 N_XI0.XI118.XI1.NET6_XI0.XI118.XI1.XI1.MM3_d
+ N_XI0.P4_XI0.XI118.XI1.XI1.MM3_g N_VDD_XI0.XI118.XI1.XI1.MM3_s
+ N_VDD_XI0.XI102.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.65e-13
+ PD=7.4e-07 PS=2.52e-06
mXI0.XI91.XI1.XI1.MM3 N_XI0.XI91.XI1.NET6_XI0.XI91.XI1.XI1.MM3_d
+ N_XI0.P3_XI0.XI91.XI1.XI1.MM3_g N_VDD_XI0.XI91.XI1.XI1.MM3_s
+ N_VDD_XI0.XI88.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.65e-13
+ PD=7.4e-07 PS=2.52e-06
mXI0.XI90.XI1.XI1.MM3 N_XI0.XI90.XI1.NET6_XI0.XI90.XI1.XI1.MM3_d
+ N_XI0.P2_XI0.XI90.XI1.XI1.MM3_g N_VDD_XI0.XI90.XI1.XI1.MM3_s
+ N_VDD_XI0.XI82.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.65e-13
+ PD=7.4e-07 PS=2.52e-06
mXI0.XI89.XI1.XI1.MM3 N_XI0.XI89.XI1.NET6_XI0.XI89.XI1.XI1.MM3_d
+ N_XI0.P1_XI0.XI89.XI1.XI1.MM3_g N_VDD_XI0.XI89.XI1.XI1.MM3_s
+ N_VDD_XI0.XI10.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.65e-13
+ PD=7.4e-07 PS=2.52e-06
mXI2.MM1 N_NET0858_XI2.MM1_d N_NET141_XI2.MM1_g N_VDD_XI2.MM1_s N_VDD_XI2.MM1_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI0.XI182.MM3 N_NET141_XI0.XI182.MM3_d N_XI0.XI182.NET39_XI0.XI182.MM3_g
+ N_XI0.XI182.NET37_XI0.XI182.MM3_s N_VDD_XI0.XI134.XI9.MM1_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.425e-12 AS=5.4375e-13 PD=1.9e-06 PS=7.25e-07
mXI0.XI168.XI1.XI0.MM1 N_XI0.XI168.NET13_XI0.XI168.XI1.XI0.MM1_d
+ N_XI0.XI168.XI1.NET6_XI0.XI168.XI1.XI0.MM1_g N_VDD_XI0.XI168.XI1.XI0.MM1_s
+ N_VDD_XI0.XI153.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI0.XI167.XI1.XI0.MM1 N_XI0.XI167.NET13_XI0.XI167.XI1.XI0.MM1_d
+ N_XI0.XI167.XI1.NET6_XI0.XI167.XI1.XI0.MM1_g N_VDD_XI0.XI167.XI1.XI0.MM1_s
+ N_VDD_XI0.XI154.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI0.XI166.XI1.XI0.MM1 N_XI0.XI166.NET13_XI0.XI166.XI1.XI0.MM1_d
+ N_XI0.XI166.XI1.NET6_XI0.XI166.XI1.XI0.MM1_g N_VDD_XI0.XI166.XI1.XI0.MM1_s
+ N_VDD_XI0.XI157.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI0.XI165.XI1.XI0.MM1 N_XI0.XI165.NET13_XI0.XI165.XI1.XI0.MM1_d
+ N_XI0.XI165.XI1.NET6_XI0.XI165.XI1.XI0.MM1_g N_VDD_XI0.XI165.XI1.XI0.MM1_s
+ N_VDD_XI0.XI156.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI0.XI159.XI1.XI0.MM1 N_XI0.XI159.NET13_XI0.XI159.XI1.XI0.MM1_d
+ N_XI0.XI159.XI1.NET6_XI0.XI159.XI1.XI0.MM1_g N_VDD_XI0.XI159.XI1.XI0.MM1_s
+ N_VDD_XI0.XI155.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI0.XI160.XI1.XI0.MM1 N_XI0.XI160.NET13_XI0.XI160.XI1.XI0.MM1_d
+ N_XI0.XI160.XI1.NET6_XI0.XI160.XI1.XI0.MM1_g N_VDD_XI0.XI160.XI1.XI0.MM1_s
+ N_VDD_XI0.XI133.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI0.XI161.XI1.XI0.MM1 N_XI0.XI161.NET13_XI0.XI161.XI1.XI0.MM1_d
+ N_XI0.XI161.XI1.NET6_XI0.XI161.XI1.XI0.MM1_g N_VDD_XI0.XI161.XI1.XI0.MM1_s
+ N_VDD_XI0.XI132.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI0.XI162.XI1.XI0.MM1 N_XI0.XI162.NET13_XI0.XI162.XI1.XI0.MM1_d
+ N_XI0.XI162.XI1.NET6_XI0.XI162.XI1.XI0.MM1_g N_VDD_XI0.XI162.XI1.XI0.MM1_s
+ N_VDD_XI0.XI131.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI0.XI121.XI1.XI0.MM1 N_XI0.XI121.NET13_XI0.XI121.XI1.XI0.MM1_d
+ N_XI0.XI121.XI1.NET6_XI0.XI121.XI1.XI0.MM1_g N_VDD_XI0.XI121.XI1.XI0.MM1_s
+ N_VDD_XI0.XI111.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI0.XI120.XI1.XI0.MM1 N_XI0.XI120.NET13_XI0.XI120.XI1.XI0.MM1_d
+ N_XI0.XI120.XI1.NET6_XI0.XI120.XI1.XI0.MM1_g N_VDD_XI0.XI120.XI1.XI0.MM1_s
+ N_VDD_XI0.XI110.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI0.XI119.XI1.XI0.MM1 N_XI0.XI119.NET13_XI0.XI119.XI1.XI0.MM1_d
+ N_XI0.XI119.XI1.NET6_XI0.XI119.XI1.XI0.MM1_g N_VDD_XI0.XI119.XI1.XI0.MM1_s
+ N_VDD_XI0.XI103.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI0.XI118.XI1.XI0.MM1 N_XI0.XI118.NET13_XI0.XI118.XI1.XI0.MM1_d
+ N_XI0.XI118.XI1.NET6_XI0.XI118.XI1.XI0.MM1_g N_VDD_XI0.XI118.XI1.XI0.MM1_s
+ N_VDD_XI0.XI102.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI0.XI91.XI1.XI0.MM1 N_XI0.XI91.NET13_XI0.XI91.XI1.XI0.MM1_d
+ N_XI0.XI91.XI1.NET6_XI0.XI91.XI1.XI0.MM1_g N_VDD_XI0.XI91.XI1.XI0.MM1_s
+ N_VDD_XI0.XI88.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI0.XI90.XI1.XI0.MM1 N_XI0.XI90.NET13_XI0.XI90.XI1.XI0.MM1_d
+ N_XI0.XI90.XI1.NET6_XI0.XI90.XI1.XI0.MM1_g N_VDD_XI0.XI90.XI1.XI0.MM1_s
+ N_VDD_XI0.XI82.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI0.XI89.XI1.XI0.MM1 N_XI0.XI89.NET13_XI0.XI89.XI1.XI0.MM1_d
+ N_XI0.XI89.XI1.NET6_XI0.XI89.XI1.XI0.MM1_g N_VDD_XI0.XI89.XI1.XI0.MM1_s
+ N_VDD_XI0.XI10.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI0.XI182.MM1 N_XI0.XI182.NET37_XI0.XI182.MM1_d N_XI0.P16_XI0.XI182.MM1_g
+ N_VDD_XI0.XI182.MM1_s N_VDD_XI0.XI134.XI9.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=5.4375e-13 AS=7.65e-13 PD=7.25e-07 PS=2.52e-06
mXI0.XI168.XI0.XI0.MM1 N_XI0.XI168.XI0.XI0.NET17_XI0.XI168.XI0.XI0.MM1_d
+ N_XI0.XI168.NET13_XI0.XI168.XI0.XI0.MM1_g N_VDD_XI0.XI168.XI0.XI0.MM1_s
+ N_VDD_XI0.XI153.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=4.125e-13 AS=7.35e-13
+ PD=5.5e-07 PS=2.48e-06
mXI0.XI167.XI0.XI0.MM1 N_XI0.XI167.XI0.XI0.NET17_XI0.XI167.XI0.XI0.MM1_d
+ N_XI0.XI167.NET13_XI0.XI167.XI0.XI0.MM1_g N_VDD_XI0.XI167.XI0.XI0.MM1_s
+ N_VDD_XI0.XI154.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=4.125e-13 AS=7.35e-13
+ PD=5.5e-07 PS=2.48e-06
mXI0.XI166.XI0.XI0.MM1 N_XI0.XI166.XI0.XI0.NET17_XI0.XI166.XI0.XI0.MM1_d
+ N_XI0.XI166.NET13_XI0.XI166.XI0.XI0.MM1_g N_VDD_XI0.XI166.XI0.XI0.MM1_s
+ N_VDD_XI0.XI157.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=4.125e-13 AS=7.35e-13
+ PD=5.5e-07 PS=2.48e-06
mXI0.XI165.XI0.XI0.MM1 N_XI0.XI165.XI0.XI0.NET17_XI0.XI165.XI0.XI0.MM1_d
+ N_XI0.XI165.NET13_XI0.XI165.XI0.XI0.MM1_g N_VDD_XI0.XI165.XI0.XI0.MM1_s
+ N_VDD_XI0.XI156.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=4.125e-13 AS=7.35e-13
+ PD=5.5e-07 PS=2.48e-06
mXI0.XI159.XI0.XI0.MM1 N_XI0.XI159.XI0.XI0.NET17_XI0.XI159.XI0.XI0.MM1_d
+ N_XI0.XI159.NET13_XI0.XI159.XI0.XI0.MM1_g N_VDD_XI0.XI159.XI0.XI0.MM1_s
+ N_VDD_XI0.XI155.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=4.125e-13 AS=7.35e-13
+ PD=5.5e-07 PS=2.48e-06
mXI0.XI160.XI0.XI0.MM1 N_XI0.XI160.XI0.XI0.NET17_XI0.XI160.XI0.XI0.MM1_d
+ N_XI0.XI160.NET13_XI0.XI160.XI0.XI0.MM1_g N_VDD_XI0.XI160.XI0.XI0.MM1_s
+ N_VDD_XI0.XI133.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=4.125e-13 AS=7.35e-13
+ PD=5.5e-07 PS=2.48e-06
mXI0.XI161.XI0.XI0.MM1 N_XI0.XI161.XI0.XI0.NET17_XI0.XI161.XI0.XI0.MM1_d
+ N_XI0.XI161.NET13_XI0.XI161.XI0.XI0.MM1_g N_VDD_XI0.XI161.XI0.XI0.MM1_s
+ N_VDD_XI0.XI132.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=4.125e-13 AS=7.35e-13
+ PD=5.5e-07 PS=2.48e-06
mXI0.XI162.XI0.XI0.MM1 N_XI0.XI162.XI0.XI0.NET17_XI0.XI162.XI0.XI0.MM1_d
+ N_XI0.XI162.NET13_XI0.XI162.XI0.XI0.MM1_g N_VDD_XI0.XI162.XI0.XI0.MM1_s
+ N_VDD_XI0.XI131.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=4.125e-13 AS=7.35e-13
+ PD=5.5e-07 PS=2.48e-06
mXI0.XI121.XI0.XI0.MM1 N_XI0.XI121.XI0.XI0.NET17_XI0.XI121.XI0.XI0.MM1_d
+ N_XI0.XI121.NET13_XI0.XI121.XI0.XI0.MM1_g N_VDD_XI0.XI121.XI0.XI0.MM1_s
+ N_VDD_XI0.XI111.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=4.125e-13 AS=7.35e-13
+ PD=5.5e-07 PS=2.48e-06
mXI0.XI120.XI0.XI0.MM1 N_XI0.XI120.XI0.XI0.NET17_XI0.XI120.XI0.XI0.MM1_d
+ N_XI0.XI120.NET13_XI0.XI120.XI0.XI0.MM1_g N_VDD_XI0.XI120.XI0.XI0.MM1_s
+ N_VDD_XI0.XI110.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=4.125e-13 AS=7.35e-13
+ PD=5.5e-07 PS=2.48e-06
mXI0.XI119.XI0.XI0.MM1 N_XI0.XI119.XI0.XI0.NET17_XI0.XI119.XI0.XI0.MM1_d
+ N_XI0.XI119.NET13_XI0.XI119.XI0.XI0.MM1_g N_VDD_XI0.XI119.XI0.XI0.MM1_s
+ N_VDD_XI0.XI103.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=4.125e-13 AS=7.35e-13
+ PD=5.5e-07 PS=2.48e-06
mXI0.XI118.XI0.XI0.MM1 N_XI0.XI118.XI0.XI0.NET17_XI0.XI118.XI0.XI0.MM1_d
+ N_XI0.XI118.NET13_XI0.XI118.XI0.XI0.MM1_g N_VDD_XI0.XI118.XI0.XI0.MM1_s
+ N_VDD_XI0.XI102.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=4.125e-13 AS=7.35e-13
+ PD=5.5e-07 PS=2.48e-06
mXI0.XI91.XI0.XI0.MM1 N_XI0.XI91.XI0.XI0.NET17_XI0.XI91.XI0.XI0.MM1_d
+ N_XI0.XI91.NET13_XI0.XI91.XI0.XI0.MM1_g N_VDD_XI0.XI91.XI0.XI0.MM1_s
+ N_VDD_XI0.XI88.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=4.125e-13 AS=7.35e-13
+ PD=5.5e-07 PS=2.48e-06
mXI0.XI90.XI0.XI0.MM1 N_XI0.XI90.XI0.XI0.NET17_XI0.XI90.XI0.XI0.MM1_d
+ N_XI0.XI90.NET13_XI0.XI90.XI0.XI0.MM1_g N_VDD_XI0.XI90.XI0.XI0.MM1_s
+ N_VDD_XI0.XI82.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=4.125e-13 AS=7.35e-13
+ PD=5.5e-07 PS=2.48e-06
mXI0.XI89.XI0.XI0.MM1 N_XI0.XI89.XI0.XI0.NET17_XI0.XI89.XI0.XI0.MM1_d
+ N_XI0.XI89.NET13_XI0.XI89.XI0.XI0.MM1_g N_VDD_XI0.XI89.XI0.XI0.MM1_s
+ N_VDD_XI0.XI10.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=4.125e-13 AS=7.35e-13
+ PD=5.5e-07 PS=2.48e-06
mXI0.XI182.XI4.MM1 N_XI0.XI182.NET39_XI0.XI182.XI4.MM1_d
+ N_XI0.NET198_XI0.XI182.XI4.MM1_g N_VDD_XI0.XI182.XI4.MM1_s
+ N_VDD_XI0.XI134.XI9.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI0.XI168.XI0.XI0.MM3 N_XI0.XI168.XI0.NET12_XI0.XI168.XI0.XI0.MM3_d
+ N_XI0.G15_XI0.XI168.XI0.XI0.MM3_g
+ N_XI0.XI168.XI0.XI0.NET17_XI0.XI168.XI0.XI0.MM3_s N_VDD_XI0.XI153.XI1.MM3_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=4.125e-13 PD=2.52e-06 PS=5.5e-07
mXI0.XI167.XI0.XI0.MM3 N_XI0.XI167.XI0.NET12_XI0.XI167.XI0.XI0.MM3_d
+ N_XI0.G14_XI0.XI167.XI0.XI0.MM3_g
+ N_XI0.XI167.XI0.XI0.NET17_XI0.XI167.XI0.XI0.MM3_s N_VDD_XI0.XI154.XI1.MM3_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=4.125e-13 PD=2.52e-06 PS=5.5e-07
mXI0.XI166.XI0.XI0.MM3 N_XI0.XI166.XI0.NET12_XI0.XI166.XI0.XI0.MM3_d
+ N_XI0.G13_XI0.XI166.XI0.XI0.MM3_g
+ N_XI0.XI166.XI0.XI0.NET17_XI0.XI166.XI0.XI0.MM3_s N_VDD_XI0.XI157.XI1.MM3_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=4.125e-13 PD=2.52e-06 PS=5.5e-07
mXI0.XI165.XI0.XI0.MM3 N_XI0.XI165.XI0.NET12_XI0.XI165.XI0.XI0.MM3_d
+ N_XI0.G12_XI0.XI165.XI0.XI0.MM3_g
+ N_XI0.XI165.XI0.XI0.NET17_XI0.XI165.XI0.XI0.MM3_s N_VDD_XI0.XI156.XI1.MM3_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=4.125e-13 PD=2.52e-06 PS=5.5e-07
mXI0.XI159.XI0.XI0.MM3 N_XI0.XI159.XI0.NET12_XI0.XI159.XI0.XI0.MM3_d
+ N_XI0.G11_XI0.XI159.XI0.XI0.MM3_g
+ N_XI0.XI159.XI0.XI0.NET17_XI0.XI159.XI0.XI0.MM3_s N_VDD_XI0.XI155.XI1.MM3_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=4.125e-13 PD=2.52e-06 PS=5.5e-07
mXI0.XI160.XI0.XI0.MM3 N_XI0.XI160.XI0.NET12_XI0.XI160.XI0.XI0.MM3_d
+ N_XI0.G10_XI0.XI160.XI0.XI0.MM3_g
+ N_XI0.XI160.XI0.XI0.NET17_XI0.XI160.XI0.XI0.MM3_s N_VDD_XI0.XI133.XI1.MM3_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=4.125e-13 PD=2.52e-06 PS=5.5e-07
mXI0.XI161.XI0.XI0.MM3 N_XI0.XI161.XI0.NET12_XI0.XI161.XI0.XI0.MM3_d
+ N_XI0.G9_XI0.XI161.XI0.XI0.MM3_g
+ N_XI0.XI161.XI0.XI0.NET17_XI0.XI161.XI0.XI0.MM3_s N_VDD_XI0.XI132.XI1.MM3_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=4.125e-13 PD=2.52e-06 PS=5.5e-07
mXI0.XI162.XI0.XI0.MM3 N_XI0.XI162.XI0.NET12_XI0.XI162.XI0.XI0.MM3_d
+ N_XI0.G8_XI0.XI162.XI0.XI0.MM3_g
+ N_XI0.XI162.XI0.XI0.NET17_XI0.XI162.XI0.XI0.MM3_s N_VDD_XI0.XI131.XI1.MM3_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=4.125e-13 PD=2.52e-06 PS=5.5e-07
mXI0.XI121.XI0.XI0.MM3 N_XI0.XI121.XI0.NET12_XI0.XI121.XI0.XI0.MM3_d
+ N_XI0.G7_XI0.XI121.XI0.XI0.MM3_g
+ N_XI0.XI121.XI0.XI0.NET17_XI0.XI121.XI0.XI0.MM3_s N_VDD_XI0.XI111.XI1.MM3_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=4.125e-13 PD=2.52e-06 PS=5.5e-07
mXI0.XI120.XI0.XI0.MM3 N_XI0.XI120.XI0.NET12_XI0.XI120.XI0.XI0.MM3_d
+ N_XI0.G6_XI0.XI120.XI0.XI0.MM3_g
+ N_XI0.XI120.XI0.XI0.NET17_XI0.XI120.XI0.XI0.MM3_s N_VDD_XI0.XI110.XI1.MM3_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=4.125e-13 PD=2.52e-06 PS=5.5e-07
mXI0.XI119.XI0.XI0.MM3 N_XI0.XI119.XI0.NET12_XI0.XI119.XI0.XI0.MM3_d
+ N_XI0.G5_XI0.XI119.XI0.XI0.MM3_g
+ N_XI0.XI119.XI0.XI0.NET17_XI0.XI119.XI0.XI0.MM3_s N_VDD_XI0.XI103.XI1.MM3_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=4.125e-13 PD=2.52e-06 PS=5.5e-07
mXI0.XI118.XI0.XI0.MM3 N_XI0.XI118.XI0.NET12_XI0.XI118.XI0.XI0.MM3_d
+ N_XI0.G4_XI0.XI118.XI0.XI0.MM3_g
+ N_XI0.XI118.XI0.XI0.NET17_XI0.XI118.XI0.XI0.MM3_s N_VDD_XI0.XI102.XI1.MM3_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=4.125e-13 PD=2.52e-06 PS=5.5e-07
mXI0.XI91.XI0.XI0.MM3 N_XI0.XI91.XI0.NET12_XI0.XI91.XI0.XI0.MM3_d
+ N_XI0.G3_XI0.XI91.XI0.XI0.MM3_g
+ N_XI0.XI91.XI0.XI0.NET17_XI0.XI91.XI0.XI0.MM3_s N_VDD_XI0.XI88.XI1.MM3_b P_18
+ L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=4.125e-13 PD=2.52e-06 PS=5.5e-07
mXI0.XI90.XI0.XI0.MM3 N_XI0.XI90.XI0.NET12_XI0.XI90.XI0.XI0.MM3_d
+ N_XI0.G2_XI0.XI90.XI0.XI0.MM3_g
+ N_XI0.XI90.XI0.XI0.NET17_XI0.XI90.XI0.XI0.MM3_s N_VDD_XI0.XI82.XI1.MM3_b P_18
+ L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=4.125e-13 PD=2.52e-06 PS=5.5e-07
mXI0.XI89.XI0.XI0.MM3 N_XI0.XI89.XI0.NET12_XI0.XI89.XI0.XI0.MM3_d
+ N_XI0.G1_XI0.XI89.XI0.XI0.MM3_g
+ N_XI0.XI89.XI0.XI0.NET17_XI0.XI89.XI0.XI0.MM3_s N_VDD_XI0.XI10.XI1.MM3_b P_18
+ L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=4.125e-13 PD=2.52e-06 PS=5.5e-07
mXI0.XI168.XI0.XI1.MM1 N_XI0.NET198_XI0.XI168.XI0.XI1.MM1_d
+ N_XI0.XI168.XI0.NET12_XI0.XI168.XI0.XI1.MM1_g N_VDD_XI0.XI168.XI0.XI1.MM1_s
+ N_VDD_XI0.XI153.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI0.XI167.XI0.XI1.MM1 N_XI0.NET288_XI0.XI167.XI0.XI1.MM1_d
+ N_XI0.XI167.XI0.NET12_XI0.XI167.XI0.XI1.MM1_g N_VDD_XI0.XI167.XI0.XI1.MM1_s
+ N_VDD_XI0.XI154.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI0.XI166.XI0.XI1.MM1 N_XI0.NET282_XI0.XI166.XI0.XI1.MM1_d
+ N_XI0.XI166.XI0.NET12_XI0.XI166.XI0.XI1.MM1_g N_VDD_XI0.XI166.XI0.XI1.MM1_s
+ N_VDD_XI0.XI157.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI0.XI165.XI0.XI1.MM1 N_XI0.NET276_XI0.XI165.XI0.XI1.MM1_d
+ N_XI0.XI165.XI0.NET12_XI0.XI165.XI0.XI1.MM1_g N_VDD_XI0.XI165.XI0.XI1.MM1_s
+ N_VDD_XI0.XI156.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI0.XI159.XI0.XI1.MM1 N_XI0.NET270_XI0.XI159.XI0.XI1.MM1_d
+ N_XI0.XI159.XI0.NET12_XI0.XI159.XI0.XI1.MM1_g N_VDD_XI0.XI159.XI0.XI1.MM1_s
+ N_VDD_XI0.XI155.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI0.XI160.XI0.XI1.MM1 N_XI0.NET246_XI0.XI160.XI0.XI1.MM1_d
+ N_XI0.XI160.XI0.NET12_XI0.XI160.XI0.XI1.MM1_g N_VDD_XI0.XI160.XI0.XI1.MM1_s
+ N_VDD_XI0.XI133.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI0.XI161.XI0.XI1.MM1 N_XI0.NET252_XI0.XI161.XI0.XI1.MM1_d
+ N_XI0.XI161.XI0.NET12_XI0.XI161.XI0.XI1.MM1_g N_VDD_XI0.XI161.XI0.XI1.MM1_s
+ N_VDD_XI0.XI132.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI0.XI162.XI0.XI1.MM1 N_XI0.NET258_XI0.XI162.XI0.XI1.MM1_d
+ N_XI0.XI162.XI0.NET12_XI0.XI162.XI0.XI1.MM1_g N_VDD_XI0.XI162.XI0.XI1.MM1_s
+ N_VDD_XI0.XI131.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI0.XI121.XI0.XI1.MM1 N_XI0.NET264_XI0.XI121.XI0.XI1.MM1_d
+ N_XI0.XI121.XI0.NET12_XI0.XI121.XI0.XI1.MM1_g N_VDD_XI0.XI121.XI0.XI1.MM1_s
+ N_VDD_XI0.XI111.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI0.XI120.XI0.XI1.MM1 N_XI0.NET204_XI0.XI120.XI0.XI1.MM1_d
+ N_XI0.XI120.XI0.NET12_XI0.XI120.XI0.XI1.MM1_g N_VDD_XI0.XI120.XI0.XI1.MM1_s
+ N_VDD_XI0.XI110.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI0.XI119.XI0.XI1.MM1 N_XI0.NET210_XI0.XI119.XI0.XI1.MM1_d
+ N_XI0.XI119.XI0.NET12_XI0.XI119.XI0.XI1.MM1_g N_VDD_XI0.XI119.XI0.XI1.MM1_s
+ N_VDD_XI0.XI103.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI0.XI118.XI0.XI1.MM1 N_XI0.NET216_XI0.XI118.XI0.XI1.MM1_d
+ N_XI0.XI118.XI0.NET12_XI0.XI118.XI0.XI1.MM1_g N_VDD_XI0.XI118.XI0.XI1.MM1_s
+ N_VDD_XI0.XI102.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI0.XI91.XI0.XI1.MM1 N_XI0.NET222_XI0.XI91.XI0.XI1.MM1_d
+ N_XI0.XI91.XI0.NET12_XI0.XI91.XI0.XI1.MM1_g N_VDD_XI0.XI91.XI0.XI1.MM1_s
+ N_VDD_XI0.XI88.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI0.XI90.XI0.XI1.MM1 N_XI0.NET228_XI0.XI90.XI0.XI1.MM1_d
+ N_XI0.XI90.XI0.NET12_XI0.XI90.XI0.XI1.MM1_g N_VDD_XI0.XI90.XI0.XI1.MM1_s
+ N_VDD_XI0.XI82.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI0.XI89.XI0.XI1.MM1 N_XI0.NET240_XI0.XI89.XI0.XI1.MM1_d
+ N_XI0.XI89.XI0.NET12_XI0.XI89.XI0.XI1.MM1_g N_VDD_XI0.XI89.XI0.XI1.MM1_s
+ N_VDD_XI0.XI10.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI18.XI18.MM1 N_NET241_XI18.XI18.MM1_d N_NET0859_XI18.XI18.MM1_g
+ N_NET508_XI18.XI18.MM1_s N_VDD_XI0.XI134.XI9.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=9.225e-13 PD=2.48e-06 PS=1.23e-06
mXI18.XI19.MM1 N_NET242_XI18.XI19.MM1_d N_NET0859_XI18.XI19.MM1_g
+ N_NET509_XI18.XI19.MM1_s N_VDD_XI0.XI153.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=9.225e-13 PD=2.48e-06 PS=1.23e-06
mXI18.XI17.MM1 N_NET243_XI18.XI17.MM1_d N_NET0859_XI18.XI17.MM1_g
+ N_NET510_XI18.XI17.MM1_s N_VDD_XI0.XI154.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=9.225e-13 PD=2.48e-06 PS=1.23e-06
mXI18.XI16.MM1 N_NET244_XI18.XI16.MM1_d N_NET0859_XI18.XI16.MM1_g
+ N_NET511_XI18.XI16.MM1_s N_VDD_XI0.XI157.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=9.225e-13 PD=2.48e-06 PS=1.23e-06
mXI18.XI21.MM1 N_NET245_XI18.XI21.MM1_d N_NET0859_XI18.XI21.MM1_g
+ N_NET512_XI18.XI21.MM1_s N_VDD_XI0.XI156.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=9.225e-13 PD=2.48e-06 PS=1.23e-06
mXI18.XI20.MM1 N_NET246_XI18.XI20.MM1_d N_NET0859_XI18.XI20.MM1_g
+ N_NET513_XI18.XI20.MM1_s N_VDD_XI0.XI155.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=9.225e-13 PD=2.48e-06 PS=1.23e-06
mXI18.XI22.MM1 N_NET247_XI18.XI22.MM1_d N_NET0859_XI18.XI22.MM1_g
+ N_NET514_XI18.XI22.MM1_s N_VDD_XI0.XI133.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=9.225e-13 PD=2.48e-06 PS=1.23e-06
mXI18.XI6.MM1 N_NET248_XI18.XI6.MM1_d N_NET0859_XI18.XI6.MM1_g
+ N_NET515_XI18.XI6.MM1_s N_VDD_XI0.XI132.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=9.225e-13 PD=2.48e-06 PS=1.23e-06
mXI18.XI5.MM1 N_NET249_XI18.XI5.MM1_d N_NET0859_XI18.XI5.MM1_g
+ N_NET516_XI18.XI5.MM1_s N_VDD_XI0.XI131.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=9.225e-13 PD=2.48e-06 PS=1.23e-06
mXI18.XI7.MM1 N_NET250_XI18.XI7.MM1_d N_NET0859_XI18.XI7.MM1_g
+ N_NET517_XI18.XI7.MM1_s N_VDD_XI0.XI111.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=9.225e-13 PD=2.48e-06 PS=1.23e-06
mXI18.XI8.MM1 N_NET251_XI18.XI8.MM1_d N_NET0859_XI18.XI8.MM1_g
+ N_NET518_XI18.XI8.MM1_s N_VDD_XI0.XI110.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=9.225e-13 PD=2.48e-06 PS=1.23e-06
mXI18.XI3.MM1 N_NET252_XI18.XI3.MM1_d N_NET0859_XI18.XI3.MM1_g
+ N_NET519_XI18.XI3.MM1_s N_VDD_XI0.XI103.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=9.225e-13 PD=2.48e-06 PS=1.23e-06
mXI18.XI4.MM1 N_NET253_XI18.XI4.MM1_d N_NET0859_XI18.XI4.MM1_g
+ N_NET520_XI18.XI4.MM1_s N_VDD_XI0.XI102.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=9.225e-13 PD=2.48e-06 PS=1.23e-06
mXI18.XI2.MM1 N_NET254_XI18.XI2.MM1_d N_NET0859_XI18.XI2.MM1_g
+ N_NET521_XI18.XI2.MM1_s N_VDD_XI0.XI88.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=9.225e-13 PD=2.48e-06 PS=1.23e-06
mXI18.XI1.MM1 N_NET255_XI18.XI1.MM1_d N_NET0859_XI18.XI1.MM1_g
+ N_NET522_XI18.XI1.MM1_s N_VDD_XI0.XI82.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=9.225e-13 PD=2.48e-06 PS=1.23e-06
mXI18.XI0.MM1 N_NET256_XI18.XI0.MM1_d N_NET0859_XI18.XI0.MM1_g
+ N_NET523_XI18.XI0.MM1_s N_VDD_XI18.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=9.225e-13 PD=2.48e-06 PS=1.23e-06
mXI18.XI18.MM0 N_MIN15_XI18.XI18.MM0_d N_XI18.XI18.NET7_XI18.XI18.MM0_g
+ N_NET508_XI18.XI18.MM0_s N_VDD_XI0.XI134.XI9.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=1.815e-12 AS=9.225e-13 PD=3.92e-06 PS=1.23e-06
mXI18.XI19.MM0 N_MIN14_XI18.XI19.MM0_d N_XI18.XI19.NET7_XI18.XI19.MM0_g
+ N_NET509_XI18.XI19.MM0_s N_VDD_XI0.XI153.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=1.815e-12 AS=9.225e-13 PD=3.92e-06 PS=1.23e-06
mXI18.XI17.MM0 N_MIN13_XI18.XI17.MM0_d N_XI18.XI17.NET7_XI18.XI17.MM0_g
+ N_NET510_XI18.XI17.MM0_s N_VDD_XI0.XI154.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=1.815e-12 AS=9.225e-13 PD=3.92e-06 PS=1.23e-06
mXI18.XI16.MM0 N_MIN12_XI18.XI16.MM0_d N_XI18.XI16.NET7_XI18.XI16.MM0_g
+ N_NET511_XI18.XI16.MM0_s N_VDD_XI0.XI157.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=1.815e-12 AS=9.225e-13 PD=3.92e-06 PS=1.23e-06
mXI18.XI21.MM0 N_MIN11_XI18.XI21.MM0_d N_XI18.XI21.NET7_XI18.XI21.MM0_g
+ N_NET512_XI18.XI21.MM0_s N_VDD_XI0.XI156.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=1.815e-12 AS=9.225e-13 PD=3.92e-06 PS=1.23e-06
mXI18.XI20.MM0 N_MIN10_XI18.XI20.MM0_d N_XI18.XI20.NET7_XI18.XI20.MM0_g
+ N_NET513_XI18.XI20.MM0_s N_VDD_XI0.XI155.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=1.815e-12 AS=9.225e-13 PD=3.92e-06 PS=1.23e-06
mXI18.XI22.MM0 N_MIN9_XI18.XI22.MM0_d N_XI18.XI22.NET7_XI18.XI22.MM0_g
+ N_NET514_XI18.XI22.MM0_s N_VDD_XI0.XI133.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=1.815e-12 AS=9.225e-13 PD=3.92e-06 PS=1.23e-06
mXI18.XI6.MM0 N_MIN8_XI18.XI6.MM0_d N_XI18.XI6.NET7_XI18.XI6.MM0_g
+ N_NET515_XI18.XI6.MM0_s N_VDD_XI0.XI132.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=1.815e-12 AS=9.225e-13 PD=3.92e-06 PS=1.23e-06
mXI18.XI5.MM0 N_MIN7_XI18.XI5.MM0_d N_XI18.XI5.NET7_XI18.XI5.MM0_g
+ N_NET516_XI18.XI5.MM0_s N_VDD_XI0.XI131.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=1.815e-12 AS=9.225e-13 PD=3.92e-06 PS=1.23e-06
mXI18.XI7.MM0 N_MIN6_XI18.XI7.MM0_d N_XI18.XI7.NET7_XI18.XI7.MM0_g
+ N_NET517_XI18.XI7.MM0_s N_VDD_XI0.XI111.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=1.815e-12 AS=9.225e-13 PD=3.92e-06 PS=1.23e-06
mXI18.XI8.MM0 N_MIN5_XI18.XI8.MM0_d N_XI18.XI8.NET7_XI18.XI8.MM0_g
+ N_NET518_XI18.XI8.MM0_s N_VDD_XI0.XI110.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=1.815e-12 AS=9.225e-13 PD=3.92e-06 PS=1.23e-06
mXI18.XI3.MM0 N_MIN4_XI18.XI3.MM0_d N_XI18.XI3.NET7_XI18.XI3.MM0_g
+ N_NET519_XI18.XI3.MM0_s N_VDD_XI0.XI103.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=1.815e-12 AS=9.225e-13 PD=3.92e-06 PS=1.23e-06
mXI18.XI4.MM0 N_MIN3_XI18.XI4.MM0_d N_XI18.XI4.NET7_XI18.XI4.MM0_g
+ N_NET520_XI18.XI4.MM0_s N_VDD_XI0.XI102.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=1.815e-12 AS=9.225e-13 PD=3.92e-06 PS=1.23e-06
mXI18.XI2.MM0 N_MIN2_XI18.XI2.MM0_d N_XI18.XI2.NET7_XI18.XI2.MM0_g
+ N_NET521_XI18.XI2.MM0_s N_VDD_XI0.XI88.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=1.815e-12 AS=9.225e-13 PD=3.92e-06 PS=1.23e-06
mXI18.XI1.MM0 N_MIN1_XI18.XI1.MM0_d N_XI18.XI1.NET7_XI18.XI1.MM0_g
+ N_NET522_XI18.XI1.MM0_s N_VDD_XI0.XI82.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=1.815e-12 AS=9.225e-13 PD=3.92e-06 PS=1.23e-06
mXI18.XI0.MM0 N_MIN0_XI18.XI0.MM0_d N_XI18.XI0.NET7_XI18.XI0.MM0_g
+ N_NET523_XI18.XI0.MM0_s N_VDD_XI18.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=1.815e-12 AS=9.225e-13 PD=3.92e-06 PS=1.23e-06
mXI18.XI18.MM5 N_XI18.XI18.NET7_XI18.XI18.MM5_d N_NET0859_XI18.XI18.MM5_g
+ N_VDD_XI18.XI18.MM5_s N_VDD_XI0.XI134.XI9.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI18.XI19.MM5 N_XI18.XI19.NET7_XI18.XI19.MM5_d N_NET0859_XI18.XI19.MM5_g
+ N_VDD_XI18.XI19.MM5_s N_VDD_XI0.XI153.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI18.XI17.MM5 N_XI18.XI17.NET7_XI18.XI17.MM5_d N_NET0859_XI18.XI17.MM5_g
+ N_VDD_XI18.XI17.MM5_s N_VDD_XI0.XI154.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI18.XI16.MM5 N_XI18.XI16.NET7_XI18.XI16.MM5_d N_NET0859_XI18.XI16.MM5_g
+ N_VDD_XI18.XI16.MM5_s N_VDD_XI0.XI157.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI18.XI21.MM5 N_XI18.XI21.NET7_XI18.XI21.MM5_d N_NET0859_XI18.XI21.MM5_g
+ N_VDD_XI18.XI21.MM5_s N_VDD_XI0.XI156.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI18.XI20.MM5 N_XI18.XI20.NET7_XI18.XI20.MM5_d N_NET0859_XI18.XI20.MM5_g
+ N_VDD_XI18.XI20.MM5_s N_VDD_XI0.XI155.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI18.XI22.MM5 N_XI18.XI22.NET7_XI18.XI22.MM5_d N_NET0859_XI18.XI22.MM5_g
+ N_VDD_XI18.XI22.MM5_s N_VDD_XI0.XI133.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI18.XI6.MM5 N_XI18.XI6.NET7_XI18.XI6.MM5_d N_NET0859_XI18.XI6.MM5_g
+ N_VDD_XI18.XI6.MM5_s N_VDD_XI0.XI132.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI18.XI5.MM5 N_XI18.XI5.NET7_XI18.XI5.MM5_d N_NET0859_XI18.XI5.MM5_g
+ N_VDD_XI18.XI5.MM5_s N_VDD_XI0.XI131.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI18.XI7.MM5 N_XI18.XI7.NET7_XI18.XI7.MM5_d N_NET0859_XI18.XI7.MM5_g
+ N_VDD_XI18.XI7.MM5_s N_VDD_XI0.XI111.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI18.XI8.MM5 N_XI18.XI8.NET7_XI18.XI8.MM5_d N_NET0859_XI18.XI8.MM5_g
+ N_VDD_XI18.XI8.MM5_s N_VDD_XI0.XI110.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI18.XI3.MM5 N_XI18.XI3.NET7_XI18.XI3.MM5_d N_NET0859_XI18.XI3.MM5_g
+ N_VDD_XI18.XI3.MM5_s N_VDD_XI0.XI103.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI18.XI4.MM5 N_XI18.XI4.NET7_XI18.XI4.MM5_d N_NET0859_XI18.XI4.MM5_g
+ N_VDD_XI18.XI4.MM5_s N_VDD_XI0.XI102.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI18.XI2.MM5 N_XI18.XI2.NET7_XI18.XI2.MM5_d N_NET0859_XI18.XI2.MM5_g
+ N_VDD_XI18.XI2.MM5_s N_VDD_XI0.XI88.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI18.XI1.MM5 N_XI18.XI1.NET7_XI18.XI1.MM5_d N_NET0859_XI18.XI1.MM5_g
+ N_VDD_XI18.XI1.MM5_s N_VDD_XI0.XI82.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI18.XI0.MM5 N_XI18.XI0.NET7_XI18.XI0.MM5_d N_NET0859_XI18.XI0.MM5_g
+ N_VDD_XI18.XI0.MM5_s N_VDD_XI18.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13
+ AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI15.MM0 N_XI15.NET40_XI15.MM0_d N_NET198_XI15.MM0_g N_VDD_XI15.MM0_s
+ N_VDD_XI15.MM0_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06
+ PS=2.48e-06
mXI15.XI16.XI1.MM3 N_XI15.XI16.NET6_XI15.XI16.XI1.MM3_d
+ N_NET198_XI15.XI16.XI1.MM3_g N_VDD_XI15.XI16.XI1.MM3_s N_VDD_XI15.MM0_b P_18
+ L=1.8e-07 W=1.5e-06 AD=4.125e-13 AS=7.35e-13 PD=5.5e-07 PS=2.48e-06
mXI15.XI16.XI1.MM1 N_XI15.XI16.NET6_XI15.XI16.XI1.MM1_d
+ N_NET508_XI15.XI16.XI1.MM1_g N_VDD_XI15.XI16.XI1.MM1_s N_VDD_XI15.MM0_b P_18
+ L=1.8e-07 W=1.5e-06 AD=4.125e-13 AS=7.65e-13 PD=5.5e-07 PS=2.52e-06
mXI15.XI16.XI0.MM1 N_NET417_XI15.XI16.XI0.MM1_d
+ N_XI15.XI16.NET6_XI15.XI16.XI0.MM1_g N_VDD_XI15.XI16.XI0.MM1_s
+ N_VDD_XI15.MM0_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06
+ PS=2.48e-06
mXI15.XI17.XI0.MM3 N_XI15.XI17.XI0.NET17_XI15.XI17.XI0.MM3_d
+ N_XI15.NET40_XI15.XI17.XI0.MM3_g N_VDD_XI15.XI17.XI0.MM3_s N_VDD_XI15.MM0_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=5.625e-13 AS=7.35e-13 PD=7.5e-07 PS=2.48e-06
mXI15.XI17.XI0.MM1 N_XI15.XI17.NET12_XI15.XI17.XI0.MM1_d
+ N_NET509_XI15.XI17.XI0.MM1_g N_XI15.XI17.XI0.NET17_XI15.XI17.XI0.MM1_s
+ N_VDD_XI15.MM0_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=5.625e-13 PD=2.52e-06
+ PS=7.5e-07
mXI15.XI17.XI1.MM1 N_NET418_XI15.XI17.XI1.MM1_d
+ N_XI15.XI17.NET12_XI15.XI17.XI1.MM1_g N_VDD_XI15.XI17.XI1.MM1_s
+ N_VDD_XI15.MM0_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06
+ PS=2.48e-06
mXI15.XI18.XI0.MM3 N_XI15.XI18.XI0.NET17_XI15.XI18.XI0.MM3_d
+ N_XI15.NET40_XI15.XI18.XI0.MM3_g N_VDD_XI15.XI18.XI0.MM3_s N_VDD_XI15.MM0_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=5.625e-13 AS=7.35e-13 PD=7.5e-07 PS=2.48e-06
mXI15.XI18.XI0.MM1 N_XI15.XI18.NET12_XI15.XI18.XI0.MM1_d
+ N_NET510_XI15.XI18.XI0.MM1_g N_XI15.XI18.XI0.NET17_XI15.XI18.XI0.MM1_s
+ N_VDD_XI15.MM0_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=5.625e-13 PD=2.52e-06
+ PS=7.5e-07
mXI15.XI18.XI1.MM1 N_NET419_XI15.XI18.XI1.MM1_d
+ N_XI15.XI18.NET12_XI15.XI18.XI1.MM1_g N_VDD_XI15.XI18.XI1.MM1_s
+ N_VDD_XI15.MM0_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06
+ PS=2.48e-06
mXI15.XI19.XI0.MM3 N_XI15.XI19.XI0.NET17_XI15.XI19.XI0.MM3_d
+ N_XI15.NET40_XI15.XI19.XI0.MM3_g N_VDD_XI15.XI19.XI0.MM3_s N_VDD_XI15.MM0_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=5.625e-13 AS=7.35e-13 PD=7.5e-07 PS=2.48e-06
mXI15.XI19.XI0.MM1 N_XI15.XI19.NET12_XI15.XI19.XI0.MM1_d
+ N_NET511_XI15.XI19.XI0.MM1_g N_XI15.XI19.XI0.NET17_XI15.XI19.XI0.MM1_s
+ N_VDD_XI15.MM0_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=5.625e-13 PD=2.52e-06
+ PS=7.5e-07
mXI15.XI19.XI1.MM1 N_NET420_XI15.XI19.XI1.MM1_d
+ N_XI15.XI19.NET12_XI15.XI19.XI1.MM1_g N_VDD_XI15.XI19.XI1.MM1_s
+ N_VDD_XI15.MM0_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06
+ PS=2.48e-06
mXI15.XI20.XI0.MM3 N_XI15.XI20.XI0.NET17_XI15.XI20.XI0.MM3_d
+ N_XI15.NET40_XI15.XI20.XI0.MM3_g N_VDD_XI15.XI20.XI0.MM3_s N_VDD_XI15.MM0_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=5.625e-13 AS=7.35e-13 PD=7.5e-07 PS=2.48e-06
mXI15.XI20.XI0.MM1 N_XI15.XI20.NET12_XI15.XI20.XI0.MM1_d
+ N_NET512_XI15.XI20.XI0.MM1_g N_XI15.XI20.XI0.NET17_XI15.XI20.XI0.MM1_s
+ N_VDD_XI15.MM0_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=5.625e-13 PD=2.52e-06
+ PS=7.5e-07
mXI15.XI20.XI1.MM1 N_NET421_XI15.XI20.XI1.MM1_d
+ N_XI15.XI20.NET12_XI15.XI20.XI1.MM1_g N_VDD_XI15.XI20.XI1.MM1_s
+ N_VDD_XI15.MM0_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06
+ PS=2.48e-06
mXI15.XI21.XI0.MM3 N_XI15.XI21.XI0.NET17_XI15.XI21.XI0.MM3_d
+ N_XI15.NET40_XI15.XI21.XI0.MM3_g N_VDD_XI15.XI21.XI0.MM3_s N_VDD_XI15.MM0_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=5.625e-13 AS=7.35e-13 PD=7.5e-07 PS=2.48e-06
mXI15.XI21.XI0.MM1 N_XI15.XI21.NET12_XI15.XI21.XI0.MM1_d
+ N_NET513_XI15.XI21.XI0.MM1_g N_XI15.XI21.XI0.NET17_XI15.XI21.XI0.MM1_s
+ N_VDD_XI15.MM0_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=5.625e-13 PD=2.52e-06
+ PS=7.5e-07
mXI15.XI21.XI1.MM1 N_NET422_XI15.XI21.XI1.MM1_d
+ N_XI15.XI21.NET12_XI15.XI21.XI1.MM1_g N_VDD_XI15.XI21.XI1.MM1_s
+ N_VDD_XI15.MM0_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06
+ PS=2.48e-06
mXI15.XI22.XI0.MM3 N_XI15.XI22.XI0.NET17_XI15.XI22.XI0.MM3_d
+ N_XI15.NET40_XI15.XI22.XI0.MM3_g N_VDD_XI15.XI22.XI0.MM3_s N_VDD_XI15.MM0_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=5.625e-13 AS=7.35e-13 PD=7.5e-07 PS=2.48e-06
mXI15.XI22.XI0.MM1 N_XI15.XI22.NET12_XI15.XI22.XI0.MM1_d
+ N_NET514_XI15.XI22.XI0.MM1_g N_XI15.XI22.XI0.NET17_XI15.XI22.XI0.MM1_s
+ N_VDD_XI15.MM0_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=5.625e-13 PD=2.52e-06
+ PS=7.5e-07
mXI15.XI22.XI1.MM1 N_NET423_XI15.XI22.XI1.MM1_d
+ N_XI15.XI22.NET12_XI15.XI22.XI1.MM1_g N_VDD_XI15.XI22.XI1.MM1_s
+ N_VDD_XI15.MM0_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06
+ PS=2.48e-06
mXI15.XI23.XI0.MM3 N_XI15.XI23.XI0.NET17_XI15.XI23.XI0.MM3_d
+ N_XI15.NET40_XI15.XI23.XI0.MM3_g N_VDD_XI15.XI23.XI0.MM3_s N_VDD_XI15.MM0_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=5.625e-13 AS=7.35e-13 PD=7.5e-07 PS=2.48e-06
mXI15.XI23.XI0.MM1 N_XI15.XI23.NET12_XI15.XI23.XI0.MM1_d
+ N_NET515_XI15.XI23.XI0.MM1_g N_XI15.XI23.XI0.NET17_XI15.XI23.XI0.MM1_s
+ N_VDD_XI15.MM0_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=5.625e-13 PD=2.52e-06
+ PS=7.5e-07
mXI15.XI23.XI1.MM1 N_NET424_XI15.XI23.XI1.MM1_d
+ N_XI15.XI23.NET12_XI15.XI23.XI1.MM1_g N_VDD_XI15.XI23.XI1.MM1_s
+ N_VDD_XI15.MM0_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06
+ PS=2.48e-06
mXI15.XI24.XI0.MM3 N_XI15.XI24.XI0.NET17_XI15.XI24.XI0.MM3_d
+ N_XI15.NET40_XI15.XI24.XI0.MM3_g N_VDD_XI15.XI24.XI0.MM3_s N_VDD_XI15.MM0_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=5.625e-13 AS=7.35e-13 PD=7.5e-07 PS=2.48e-06
mXI15.XI24.XI0.MM1 N_XI15.XI24.NET12_XI15.XI24.XI0.MM1_d
+ N_NET516_XI15.XI24.XI0.MM1_g N_XI15.XI24.XI0.NET17_XI15.XI24.XI0.MM1_s
+ N_VDD_XI15.MM0_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=5.625e-13 PD=2.52e-06
+ PS=7.5e-07
mXI15.XI24.XI1.MM1 N_NET425_XI15.XI24.XI1.MM1_d
+ N_XI15.XI24.NET12_XI15.XI24.XI1.MM1_g N_VDD_XI15.XI24.XI1.MM1_s
+ N_VDD_XI15.MM0_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06
+ PS=2.48e-06
mXI15.XI25.XI0.MM3 N_XI15.XI25.XI0.NET17_XI15.XI25.XI0.MM3_d
+ N_XI15.NET40_XI15.XI25.XI0.MM3_g N_VDD_XI15.XI25.XI0.MM3_s N_VDD_XI15.MM0_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=5.625e-13 AS=7.35e-13 PD=7.5e-07 PS=2.48e-06
mXI15.XI25.XI0.MM1 N_XI15.XI25.NET12_XI15.XI25.XI0.MM1_d
+ N_NET517_XI15.XI25.XI0.MM1_g N_XI15.XI25.XI0.NET17_XI15.XI25.XI0.MM1_s
+ N_VDD_XI15.MM0_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=5.625e-13 PD=2.52e-06
+ PS=7.5e-07
mXI15.XI25.XI1.MM1 N_NET426_XI15.XI25.XI1.MM1_d
+ N_XI15.XI25.NET12_XI15.XI25.XI1.MM1_g N_VDD_XI15.XI25.XI1.MM1_s
+ N_VDD_XI15.MM0_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06
+ PS=2.48e-06
mXI15.XI26.XI0.MM3 N_XI15.XI26.XI0.NET17_XI15.XI26.XI0.MM3_d
+ N_XI15.NET40_XI15.XI26.XI0.MM3_g N_VDD_XI15.XI26.XI0.MM3_s N_VDD_XI15.MM0_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=5.625e-13 AS=7.35e-13 PD=7.5e-07 PS=2.48e-06
mXI15.XI26.XI0.MM1 N_XI15.XI26.NET12_XI15.XI26.XI0.MM1_d
+ N_NET518_XI15.XI26.XI0.MM1_g N_XI15.XI26.XI0.NET17_XI15.XI26.XI0.MM1_s
+ N_VDD_XI15.MM0_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=5.625e-13 PD=2.52e-06
+ PS=7.5e-07
mXI15.XI26.XI1.MM1 N_NET427_XI15.XI26.XI1.MM1_d
+ N_XI15.XI26.NET12_XI15.XI26.XI1.MM1_g N_VDD_XI15.XI26.XI1.MM1_s
+ N_VDD_XI15.MM0_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06
+ PS=2.48e-06
mXI15.XI27.XI0.MM3 N_XI15.XI27.XI0.NET17_XI15.XI27.XI0.MM3_d
+ N_XI15.NET40_XI15.XI27.XI0.MM3_g N_VDD_XI15.XI27.XI0.MM3_s N_VDD_XI15.MM0_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=5.625e-13 AS=7.35e-13 PD=7.5e-07 PS=2.48e-06
mXI15.XI27.XI0.MM1 N_XI15.XI27.NET12_XI15.XI27.XI0.MM1_d
+ N_NET519_XI15.XI27.XI0.MM1_g N_XI15.XI27.XI0.NET17_XI15.XI27.XI0.MM1_s
+ N_VDD_XI15.MM0_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=5.625e-13 PD=2.52e-06
+ PS=7.5e-07
mXI15.XI27.XI1.MM1 N_NET428_XI15.XI27.XI1.MM1_d
+ N_XI15.XI27.NET12_XI15.XI27.XI1.MM1_g N_VDD_XI15.XI27.XI1.MM1_s
+ N_VDD_XI15.MM0_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06
+ PS=2.48e-06
mXI15.XI28.XI0.MM3 N_XI15.XI28.XI0.NET17_XI15.XI28.XI0.MM3_d
+ N_XI15.NET40_XI15.XI28.XI0.MM3_g N_VDD_XI15.XI28.XI0.MM3_s N_VDD_XI15.MM0_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=5.625e-13 AS=7.35e-13 PD=7.5e-07 PS=2.48e-06
mXI15.XI28.XI0.MM1 N_XI15.XI28.NET12_XI15.XI28.XI0.MM1_d
+ N_NET520_XI15.XI28.XI0.MM1_g N_XI15.XI28.XI0.NET17_XI15.XI28.XI0.MM1_s
+ N_VDD_XI15.MM0_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=5.625e-13 PD=2.52e-06
+ PS=7.5e-07
mXI15.XI28.XI1.MM1 N_NET429_XI15.XI28.XI1.MM1_d
+ N_XI15.XI28.NET12_XI15.XI28.XI1.MM1_g N_VDD_XI15.XI28.XI1.MM1_s
+ N_VDD_XI15.MM0_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06
+ PS=2.48e-06
mXI15.XI29.XI0.MM3 N_XI15.XI29.XI0.NET17_XI15.XI29.XI0.MM3_d
+ N_XI15.NET40_XI15.XI29.XI0.MM3_g N_VDD_XI15.XI29.XI0.MM3_s N_VDD_XI15.MM0_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=5.625e-13 AS=7.35e-13 PD=7.5e-07 PS=2.48e-06
mXI15.XI29.XI0.MM1 N_XI15.XI29.NET12_XI15.XI29.XI0.MM1_d
+ N_NET521_XI15.XI29.XI0.MM1_g N_XI15.XI29.XI0.NET17_XI15.XI29.XI0.MM1_s
+ N_VDD_XI15.MM0_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=5.625e-13 PD=2.52e-06
+ PS=7.5e-07
mXI15.XI29.XI1.MM1 N_NET430_XI15.XI29.XI1.MM1_d
+ N_XI15.XI29.NET12_XI15.XI29.XI1.MM1_g N_VDD_XI15.XI29.XI1.MM1_s
+ N_VDD_XI15.MM0_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06
+ PS=2.48e-06
mXI15.XI30.XI0.MM3 N_XI15.XI30.XI0.NET17_XI15.XI30.XI0.MM3_d
+ N_XI15.NET40_XI15.XI30.XI0.MM3_g N_VDD_XI15.XI30.XI0.MM3_s N_VDD_XI15.MM0_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=5.625e-13 AS=7.35e-13 PD=7.5e-07 PS=2.48e-06
mXI15.XI30.XI0.MM1 N_XI15.XI30.NET12_XI15.XI30.XI0.MM1_d
+ N_NET522_XI15.XI30.XI0.MM1_g N_XI15.XI30.XI0.NET17_XI15.XI30.XI0.MM1_s
+ N_VDD_XI15.MM0_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=5.625e-13 PD=2.52e-06
+ PS=7.5e-07
mXI15.XI30.XI1.MM1 N_NET431_XI15.XI30.XI1.MM1_d
+ N_XI15.XI30.NET12_XI15.XI30.XI1.MM1_g N_VDD_XI15.XI30.XI1.MM1_s
+ N_VDD_XI15.MM0_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06
+ PS=2.48e-06
mXI15.XI31.XI0.MM3 N_XI15.XI31.XI0.NET17_XI15.XI31.XI0.MM3_d
+ N_XI15.NET40_XI15.XI31.XI0.MM3_g N_VDD_XI15.XI31.XI0.MM3_s N_VDD_XI15.MM0_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=5.625e-13 AS=7.35e-13 PD=7.5e-07 PS=2.48e-06
mXI15.XI31.XI0.MM1 N_XI15.XI31.NET12_XI15.XI31.XI0.MM1_d
+ N_NET523_XI15.XI31.XI0.MM1_g N_XI15.XI31.XI0.NET17_XI15.XI31.XI0.MM1_s
+ N_VDD_XI15.MM0_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=5.625e-13 PD=2.52e-06
+ PS=7.5e-07
mXI15.XI31.XI1.MM1 N_NET432_XI15.XI31.XI1.MM1_d
+ N_XI15.XI31.NET12_XI15.XI31.XI1.MM1_g N_VDD_XI15.XI31.XI1.MM1_s
+ N_VDD_XI15.MM0_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06
+ PS=2.48e-06
mXI12.XI30.XI0.MM1 N_XI12.XI30.NET0180_XI12.XI30.XI0.MM1_d
+ N_NET222_XI12.XI30.XI0.MM1_g N_VDD_XI12.XI30.XI0.MM1_s
+ N_VDD_XI12.XI30.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI12.XI29.XI0.MM1 N_XI12.XI29.NET0180_XI12.XI29.XI0.MM1_d
+ N_NET222_XI12.XI29.XI0.MM1_g N_VDD_XI12.XI29.XI0.MM1_s
+ N_VDD_XI12.XI29.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI12.XI31.XI0.MM1 N_XI12.XI31.NET0180_XI12.XI31.XI0.MM1_d
+ N_NET222_XI12.XI31.XI0.MM1_g N_VDD_XI12.XI31.XI0.MM1_s
+ N_VDD_XI12.XI31.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI12.XI28.XI0.MM1 N_XI12.XI28.NET0180_XI12.XI28.XI0.MM1_d
+ N_NET222_XI12.XI28.XI0.MM1_g N_VDD_XI12.XI28.XI0.MM1_s
+ N_VDD_XI12.XI28.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI12.XI25.XI0.MM1 N_XI12.XI25.NET0180_XI12.XI25.XI0.MM1_d
+ N_NET222_XI12.XI25.XI0.MM1_g N_VDD_XI12.XI25.XI0.MM1_s
+ N_VDD_XI12.XI25.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI12.XI26.XI0.MM1 N_XI12.XI26.NET0180_XI12.XI26.XI0.MM1_d
+ N_NET222_XI12.XI26.XI0.MM1_g N_VDD_XI12.XI26.XI0.MM1_s
+ N_VDD_XI12.XI26.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI12.XI24.XI0.MM1 N_XI12.XI24.NET0180_XI12.XI24.XI0.MM1_d
+ N_NET222_XI12.XI24.XI0.MM1_g N_VDD_XI12.XI24.XI0.MM1_s
+ N_VDD_XI12.XI24.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI12.XI27.XI0.MM1 N_XI12.XI27.NET0180_XI12.XI27.XI0.MM1_d
+ N_NET222_XI12.XI27.XI0.MM1_g N_VDD_XI12.XI27.XI0.MM1_s
+ N_VDD_XI12.XI27.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI12.XI22.XI0.MM1 N_XI12.XI22.NET0180_XI12.XI22.XI0.MM1_d
+ N_NET222_XI12.XI22.XI0.MM1_g N_VDD_XI12.XI22.XI0.MM1_s
+ N_VDD_XI12.XI22.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI12.XI21.XI0.MM1 N_XI12.XI21.NET0180_XI12.XI21.XI0.MM1_d
+ N_NET222_XI12.XI21.XI0.MM1_g N_VDD_XI12.XI21.XI0.MM1_s
+ N_VDD_XI12.XI21.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI12.XI23.XI0.MM1 N_XI12.XI23.NET0180_XI12.XI23.XI0.MM1_d
+ N_NET222_XI12.XI23.XI0.MM1_g N_VDD_XI12.XI23.XI0.MM1_s
+ N_VDD_XI12.XI23.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI12.XI19.XI0.MM1 N_XI12.XI19.NET0180_XI12.XI19.XI0.MM1_d
+ N_NET222_XI12.XI19.XI0.MM1_g N_VDD_XI12.XI19.XI0.MM1_s
+ N_VDD_XI12.XI19.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI12.XI20.XI0.MM1 N_XI12.XI20.NET0180_XI12.XI20.XI0.MM1_d
+ N_NET222_XI12.XI20.XI0.MM1_g N_VDD_XI12.XI20.XI0.MM1_s
+ N_VDD_XI12.XI20.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI12.XI18.XI0.MM1 N_XI12.XI18.NET0180_XI12.XI18.XI0.MM1_d
+ N_NET222_XI12.XI18.XI0.MM1_g N_VDD_XI12.XI18.XI0.MM1_s
+ N_VDD_XI12.XI18.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI12.XI17.XI0.MM1 N_XI12.XI17.NET0180_XI12.XI17.XI0.MM1_d
+ N_NET222_XI12.XI17.XI0.MM1_g N_VDD_XI12.XI17.XI0.MM1_s
+ N_VDD_XI12.XI17.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI12.XI0.XI0.MM1 N_XI12.XI0.NET0180_XI12.XI0.XI0.MM1_d
+ N_NET222_XI12.XI0.XI0.MM1_g N_VDD_XI12.XI0.XI0.MM1_s N_VDD_XI12.XI0.XI0.MM1_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI12.XI30.XI1.MM1 N_XI12.XI30.NET35_XI12.XI30.XI1.MM1_d
+ N_XI12.XI30.NET0180_XI12.XI30.XI1.MM1_g N_VDD_XI12.XI30.XI1.MM1_s
+ N_VDD_XI12.XI30.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI12.XI29.XI1.MM1 N_XI12.XI29.NET35_XI12.XI29.XI1.MM1_d
+ N_XI12.XI29.NET0180_XI12.XI29.XI1.MM1_g N_VDD_XI12.XI29.XI1.MM1_s
+ N_VDD_XI12.XI29.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI12.XI31.XI1.MM1 N_XI12.XI31.NET35_XI12.XI31.XI1.MM1_d
+ N_XI12.XI31.NET0180_XI12.XI31.XI1.MM1_g N_VDD_XI12.XI31.XI1.MM1_s
+ N_VDD_XI12.XI31.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI12.XI28.XI1.MM1 N_XI12.XI28.NET35_XI12.XI28.XI1.MM1_d
+ N_XI12.XI28.NET0180_XI12.XI28.XI1.MM1_g N_VDD_XI12.XI28.XI1.MM1_s
+ N_VDD_XI12.XI28.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI12.XI25.XI1.MM1 N_XI12.XI25.NET35_XI12.XI25.XI1.MM1_d
+ N_XI12.XI25.NET0180_XI12.XI25.XI1.MM1_g N_VDD_XI12.XI25.XI1.MM1_s
+ N_VDD_XI12.XI25.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI12.XI26.XI1.MM1 N_XI12.XI26.NET35_XI12.XI26.XI1.MM1_d
+ N_XI12.XI26.NET0180_XI12.XI26.XI1.MM1_g N_VDD_XI12.XI26.XI1.MM1_s
+ N_VDD_XI12.XI26.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI12.XI24.XI1.MM1 N_XI12.XI24.NET35_XI12.XI24.XI1.MM1_d
+ N_XI12.XI24.NET0180_XI12.XI24.XI1.MM1_g N_VDD_XI12.XI24.XI1.MM1_s
+ N_VDD_XI12.XI24.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI12.XI27.XI1.MM1 N_XI12.XI27.NET35_XI12.XI27.XI1.MM1_d
+ N_XI12.XI27.NET0180_XI12.XI27.XI1.MM1_g N_VDD_XI12.XI27.XI1.MM1_s
+ N_VDD_XI12.XI27.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI12.XI22.XI1.MM1 N_XI12.XI22.NET35_XI12.XI22.XI1.MM1_d
+ N_XI12.XI22.NET0180_XI12.XI22.XI1.MM1_g N_VDD_XI12.XI22.XI1.MM1_s
+ N_VDD_XI12.XI22.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI12.XI21.XI1.MM1 N_XI12.XI21.NET35_XI12.XI21.XI1.MM1_d
+ N_XI12.XI21.NET0180_XI12.XI21.XI1.MM1_g N_VDD_XI12.XI21.XI1.MM1_s
+ N_VDD_XI12.XI21.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI12.XI23.XI1.MM1 N_XI12.XI23.NET35_XI12.XI23.XI1.MM1_d
+ N_XI12.XI23.NET0180_XI12.XI23.XI1.MM1_g N_VDD_XI12.XI23.XI1.MM1_s
+ N_VDD_XI12.XI23.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI12.XI19.XI1.MM1 N_XI12.XI19.NET35_XI12.XI19.XI1.MM1_d
+ N_XI12.XI19.NET0180_XI12.XI19.XI1.MM1_g N_VDD_XI12.XI19.XI1.MM1_s
+ N_VDD_XI12.XI19.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI12.XI20.XI1.MM1 N_XI12.XI20.NET35_XI12.XI20.XI1.MM1_d
+ N_XI12.XI20.NET0180_XI12.XI20.XI1.MM1_g N_VDD_XI12.XI20.XI1.MM1_s
+ N_VDD_XI12.XI20.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI12.XI18.XI1.MM1 N_XI12.XI18.NET35_XI12.XI18.XI1.MM1_d
+ N_XI12.XI18.NET0180_XI12.XI18.XI1.MM1_g N_VDD_XI12.XI18.XI1.MM1_s
+ N_VDD_XI12.XI18.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI12.XI17.XI1.MM1 N_XI12.XI17.NET35_XI12.XI17.XI1.MM1_d
+ N_XI12.XI17.NET0180_XI12.XI17.XI1.MM1_g N_VDD_XI12.XI17.XI1.MM1_s
+ N_VDD_XI12.XI17.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI12.XI0.XI1.MM1 N_XI12.XI0.NET35_XI12.XI0.XI1.MM1_d
+ N_XI12.XI0.NET0180_XI12.XI0.XI1.MM1_g N_VDD_XI12.XI0.XI1.MM1_s
+ N_VDD_XI12.XI0.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI12.XI30.MM25 N_XI12.XI30.CLKB_XI12.XI30.MM25_d
+ N_XI12.XI30.NET35_XI12.XI30.MM25_g N_VDD_XI12.XI30.MM25_s
+ N_VDD_XI12.XI30.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI12.XI29.MM25 N_XI12.XI29.CLKB_XI12.XI29.MM25_d
+ N_XI12.XI29.NET35_XI12.XI29.MM25_g N_VDD_XI12.XI29.MM25_s
+ N_VDD_XI12.XI29.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI12.XI31.MM25 N_XI12.XI31.CLKB_XI12.XI31.MM25_d
+ N_XI12.XI31.NET35_XI12.XI31.MM25_g N_VDD_XI12.XI31.MM25_s
+ N_VDD_XI12.XI31.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI12.XI28.MM25 N_XI12.XI28.CLKB_XI12.XI28.MM25_d
+ N_XI12.XI28.NET35_XI12.XI28.MM25_g N_VDD_XI12.XI28.MM25_s
+ N_VDD_XI12.XI28.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI12.XI25.MM25 N_XI12.XI25.CLKB_XI12.XI25.MM25_d
+ N_XI12.XI25.NET35_XI12.XI25.MM25_g N_VDD_XI12.XI25.MM25_s
+ N_VDD_XI12.XI25.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI12.XI26.MM25 N_XI12.XI26.CLKB_XI12.XI26.MM25_d
+ N_XI12.XI26.NET35_XI12.XI26.MM25_g N_VDD_XI12.XI26.MM25_s
+ N_VDD_XI12.XI26.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI12.XI24.MM25 N_XI12.XI24.CLKB_XI12.XI24.MM25_d
+ N_XI12.XI24.NET35_XI12.XI24.MM25_g N_VDD_XI12.XI24.MM25_s
+ N_VDD_XI12.XI24.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI12.XI27.MM25 N_XI12.XI27.CLKB_XI12.XI27.MM25_d
+ N_XI12.XI27.NET35_XI12.XI27.MM25_g N_VDD_XI12.XI27.MM25_s
+ N_VDD_XI12.XI27.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI12.XI22.MM25 N_XI12.XI22.CLKB_XI12.XI22.MM25_d
+ N_XI12.XI22.NET35_XI12.XI22.MM25_g N_VDD_XI12.XI22.MM25_s
+ N_VDD_XI12.XI22.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI12.XI21.MM25 N_XI12.XI21.CLKB_XI12.XI21.MM25_d
+ N_XI12.XI21.NET35_XI12.XI21.MM25_g N_VDD_XI12.XI21.MM25_s
+ N_VDD_XI12.XI21.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI12.XI23.MM25 N_XI12.XI23.CLKB_XI12.XI23.MM25_d
+ N_XI12.XI23.NET35_XI12.XI23.MM25_g N_VDD_XI12.XI23.MM25_s
+ N_VDD_XI12.XI23.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI12.XI19.MM25 N_XI12.XI19.CLKB_XI12.XI19.MM25_d
+ N_XI12.XI19.NET35_XI12.XI19.MM25_g N_VDD_XI12.XI19.MM25_s
+ N_VDD_XI12.XI19.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI12.XI20.MM25 N_XI12.XI20.CLKB_XI12.XI20.MM25_d
+ N_XI12.XI20.NET35_XI12.XI20.MM25_g N_VDD_XI12.XI20.MM25_s
+ N_VDD_XI12.XI20.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI12.XI18.MM25 N_XI12.XI18.CLKB_XI12.XI18.MM25_d
+ N_XI12.XI18.NET35_XI12.XI18.MM25_g N_VDD_XI12.XI18.MM25_s
+ N_VDD_XI12.XI18.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI12.XI17.MM25 N_XI12.XI17.CLKB_XI12.XI17.MM25_d
+ N_XI12.XI17.NET35_XI12.XI17.MM25_g N_VDD_XI12.XI17.MM25_s
+ N_VDD_XI12.XI17.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI12.XI0.MM25 N_XI12.XI0.CLKB_XI12.XI0.MM25_d N_XI12.XI0.NET35_XI12.XI0.MM25_g
+ N_VDD_XI12.XI0.MM25_s N_VDD_XI12.XI0.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI12.XI30.MM20 N_XI12.XI30.NET27_XI12.XI30.MM20_d N_NET417_XI12.XI30.MM20_g
+ N_VDD_XI12.XI30.MM20_s N_VDD_XI12.XI30.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI12.XI29.MM20 N_XI12.XI29.NET27_XI12.XI29.MM20_d N_NET418_XI12.XI29.MM20_g
+ N_VDD_XI12.XI29.MM20_s N_VDD_XI12.XI29.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI12.XI31.MM20 N_XI12.XI31.NET27_XI12.XI31.MM20_d N_NET419_XI12.XI31.MM20_g
+ N_VDD_XI12.XI31.MM20_s N_VDD_XI12.XI31.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI12.XI28.MM20 N_XI12.XI28.NET27_XI12.XI28.MM20_d N_NET420_XI12.XI28.MM20_g
+ N_VDD_XI12.XI28.MM20_s N_VDD_XI12.XI28.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI12.XI25.MM20 N_XI12.XI25.NET27_XI12.XI25.MM20_d N_NET421_XI12.XI25.MM20_g
+ N_VDD_XI12.XI25.MM20_s N_VDD_XI12.XI25.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI12.XI26.MM20 N_XI12.XI26.NET27_XI12.XI26.MM20_d N_NET422_XI12.XI26.MM20_g
+ N_VDD_XI12.XI26.MM20_s N_VDD_XI12.XI26.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI12.XI24.MM20 N_XI12.XI24.NET27_XI12.XI24.MM20_d N_NET423_XI12.XI24.MM20_g
+ N_VDD_XI12.XI24.MM20_s N_VDD_XI12.XI24.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI12.XI27.MM20 N_XI12.XI27.NET27_XI12.XI27.MM20_d N_NET424_XI12.XI27.MM20_g
+ N_VDD_XI12.XI27.MM20_s N_VDD_XI12.XI27.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI12.XI22.MM20 N_XI12.XI22.NET27_XI12.XI22.MM20_d N_NET425_XI12.XI22.MM20_g
+ N_VDD_XI12.XI22.MM20_s N_VDD_XI12.XI22.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI12.XI21.MM20 N_XI12.XI21.NET27_XI12.XI21.MM20_d N_NET426_XI12.XI21.MM20_g
+ N_VDD_XI12.XI21.MM20_s N_VDD_XI12.XI21.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI12.XI23.MM20 N_XI12.XI23.NET27_XI12.XI23.MM20_d N_NET427_XI12.XI23.MM20_g
+ N_VDD_XI12.XI23.MM20_s N_VDD_XI12.XI23.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI12.XI19.MM20 N_XI12.XI19.NET27_XI12.XI19.MM20_d N_NET428_XI12.XI19.MM20_g
+ N_VDD_XI12.XI19.MM20_s N_VDD_XI12.XI19.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI12.XI20.MM20 N_XI12.XI20.NET27_XI12.XI20.MM20_d N_NET429_XI12.XI20.MM20_g
+ N_VDD_XI12.XI20.MM20_s N_VDD_XI12.XI20.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI12.XI18.MM20 N_XI12.XI18.NET27_XI12.XI18.MM20_d N_NET430_XI12.XI18.MM20_g
+ N_VDD_XI12.XI18.MM20_s N_VDD_XI12.XI18.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI12.XI17.MM20 N_XI12.XI17.NET27_XI12.XI17.MM20_d N_NET431_XI12.XI17.MM20_g
+ N_VDD_XI12.XI17.MM20_s N_VDD_XI12.XI17.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI12.XI0.MM20 N_XI12.XI0.NET27_XI12.XI0.MM20_d N_NET432_XI12.XI0.MM20_g
+ N_VDD_XI12.XI0.MM20_s N_VDD_XI12.XI0.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI12.XI30.MM17 N_XI12.XI30.NET31_XI12.XI30.MM17_d
+ N_XI12.XI30.NET27_XI12.XI30.MM17_g N_VDD_XI12.XI30.MM17_s
+ N_VDD_XI12.XI30.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI12.XI29.MM17 N_XI12.XI29.NET31_XI12.XI29.MM17_d
+ N_XI12.XI29.NET27_XI12.XI29.MM17_g N_VDD_XI12.XI29.MM17_s
+ N_VDD_XI12.XI29.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI12.XI31.MM17 N_XI12.XI31.NET31_XI12.XI31.MM17_d
+ N_XI12.XI31.NET27_XI12.XI31.MM17_g N_VDD_XI12.XI31.MM17_s
+ N_VDD_XI12.XI31.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI12.XI28.MM17 N_XI12.XI28.NET31_XI12.XI28.MM17_d
+ N_XI12.XI28.NET27_XI12.XI28.MM17_g N_VDD_XI12.XI28.MM17_s
+ N_VDD_XI12.XI28.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI12.XI25.MM17 N_XI12.XI25.NET31_XI12.XI25.MM17_d
+ N_XI12.XI25.NET27_XI12.XI25.MM17_g N_VDD_XI12.XI25.MM17_s
+ N_VDD_XI12.XI25.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI12.XI26.MM17 N_XI12.XI26.NET31_XI12.XI26.MM17_d
+ N_XI12.XI26.NET27_XI12.XI26.MM17_g N_VDD_XI12.XI26.MM17_s
+ N_VDD_XI12.XI26.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI12.XI24.MM17 N_XI12.XI24.NET31_XI12.XI24.MM17_d
+ N_XI12.XI24.NET27_XI12.XI24.MM17_g N_VDD_XI12.XI24.MM17_s
+ N_VDD_XI12.XI24.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI12.XI27.MM17 N_XI12.XI27.NET31_XI12.XI27.MM17_d
+ N_XI12.XI27.NET27_XI12.XI27.MM17_g N_VDD_XI12.XI27.MM17_s
+ N_VDD_XI12.XI27.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI12.XI22.MM17 N_XI12.XI22.NET31_XI12.XI22.MM17_d
+ N_XI12.XI22.NET27_XI12.XI22.MM17_g N_VDD_XI12.XI22.MM17_s
+ N_VDD_XI12.XI22.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI12.XI21.MM17 N_XI12.XI21.NET31_XI12.XI21.MM17_d
+ N_XI12.XI21.NET27_XI12.XI21.MM17_g N_VDD_XI12.XI21.MM17_s
+ N_VDD_XI12.XI21.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI12.XI23.MM17 N_XI12.XI23.NET31_XI12.XI23.MM17_d
+ N_XI12.XI23.NET27_XI12.XI23.MM17_g N_VDD_XI12.XI23.MM17_s
+ N_VDD_XI12.XI23.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI12.XI19.MM17 N_XI12.XI19.NET31_XI12.XI19.MM17_d
+ N_XI12.XI19.NET27_XI12.XI19.MM17_g N_VDD_XI12.XI19.MM17_s
+ N_VDD_XI12.XI19.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI12.XI20.MM17 N_XI12.XI20.NET31_XI12.XI20.MM17_d
+ N_XI12.XI20.NET27_XI12.XI20.MM17_g N_VDD_XI12.XI20.MM17_s
+ N_VDD_XI12.XI20.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI12.XI18.MM17 N_XI12.XI18.NET31_XI12.XI18.MM17_d
+ N_XI12.XI18.NET27_XI12.XI18.MM17_g N_VDD_XI12.XI18.MM17_s
+ N_VDD_XI12.XI18.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI12.XI17.MM17 N_XI12.XI17.NET31_XI12.XI17.MM17_d
+ N_XI12.XI17.NET27_XI12.XI17.MM17_g N_VDD_XI12.XI17.MM17_s
+ N_VDD_XI12.XI17.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI12.XI0.MM17 N_XI12.XI0.NET31_XI12.XI0.MM17_d N_XI12.XI0.NET27_XI12.XI0.MM17_g
+ N_VDD_XI12.XI0.MM17_s N_VDD_XI12.XI0.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI12.XI30.MM27 N_XI12.XI30.NET31_XI12.XI30.MM27_d
+ N_XI12.XI30.NET35_XI12.XI30.MM27_g N_XI12.XI30.NET58_XI12.XI30.MM27_s
+ N_VDD_XI12.XI30.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=1.125e-12 AS=9.375e-13
+ PD=3e-06 PS=2.75e-06
mXI12.XI29.MM27 N_XI12.XI29.NET31_XI12.XI29.MM27_d
+ N_XI12.XI29.NET35_XI12.XI29.MM27_g N_XI12.XI29.NET58_XI12.XI29.MM27_s
+ N_VDD_XI12.XI29.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=1.125e-12 AS=9.375e-13
+ PD=3e-06 PS=2.75e-06
mXI12.XI31.MM27 N_XI12.XI31.NET31_XI12.XI31.MM27_d
+ N_XI12.XI31.NET35_XI12.XI31.MM27_g N_XI12.XI31.NET58_XI12.XI31.MM27_s
+ N_VDD_XI12.XI31.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=1.125e-12 AS=9.375e-13
+ PD=3e-06 PS=2.75e-06
mXI12.XI28.MM27 N_XI12.XI28.NET31_XI12.XI28.MM27_d
+ N_XI12.XI28.NET35_XI12.XI28.MM27_g N_XI12.XI28.NET58_XI12.XI28.MM27_s
+ N_VDD_XI12.XI28.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=1.125e-12 AS=9.375e-13
+ PD=3e-06 PS=2.75e-06
mXI12.XI25.MM27 N_XI12.XI25.NET31_XI12.XI25.MM27_d
+ N_XI12.XI25.NET35_XI12.XI25.MM27_g N_XI12.XI25.NET58_XI12.XI25.MM27_s
+ N_VDD_XI12.XI25.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=1.125e-12 AS=9.375e-13
+ PD=3e-06 PS=2.75e-06
mXI12.XI26.MM27 N_XI12.XI26.NET31_XI12.XI26.MM27_d
+ N_XI12.XI26.NET35_XI12.XI26.MM27_g N_XI12.XI26.NET58_XI12.XI26.MM27_s
+ N_VDD_XI12.XI26.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=1.125e-12 AS=9.375e-13
+ PD=3e-06 PS=2.75e-06
mXI12.XI24.MM27 N_XI12.XI24.NET31_XI12.XI24.MM27_d
+ N_XI12.XI24.NET35_XI12.XI24.MM27_g N_XI12.XI24.NET58_XI12.XI24.MM27_s
+ N_VDD_XI12.XI24.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=1.125e-12 AS=9.375e-13
+ PD=3e-06 PS=2.75e-06
mXI12.XI27.MM27 N_XI12.XI27.NET31_XI12.XI27.MM27_d
+ N_XI12.XI27.NET35_XI12.XI27.MM27_g N_XI12.XI27.NET58_XI12.XI27.MM27_s
+ N_VDD_XI12.XI27.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=1.125e-12 AS=9.375e-13
+ PD=3e-06 PS=2.75e-06
mXI12.XI22.MM27 N_XI12.XI22.NET31_XI12.XI22.MM27_d
+ N_XI12.XI22.NET35_XI12.XI22.MM27_g N_XI12.XI22.NET58_XI12.XI22.MM27_s
+ N_VDD_XI12.XI22.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=1.125e-12 AS=9.375e-13
+ PD=3e-06 PS=2.75e-06
mXI12.XI21.MM27 N_XI12.XI21.NET31_XI12.XI21.MM27_d
+ N_XI12.XI21.NET35_XI12.XI21.MM27_g N_XI12.XI21.NET58_XI12.XI21.MM27_s
+ N_VDD_XI12.XI21.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=1.125e-12 AS=9.375e-13
+ PD=3e-06 PS=2.75e-06
mXI12.XI23.MM27 N_XI12.XI23.NET31_XI12.XI23.MM27_d
+ N_XI12.XI23.NET35_XI12.XI23.MM27_g N_XI12.XI23.NET58_XI12.XI23.MM27_s
+ N_VDD_XI12.XI23.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=1.125e-12 AS=9.375e-13
+ PD=3e-06 PS=2.75e-06
mXI12.XI19.MM27 N_XI12.XI19.NET31_XI12.XI19.MM27_d
+ N_XI12.XI19.NET35_XI12.XI19.MM27_g N_XI12.XI19.NET58_XI12.XI19.MM27_s
+ N_VDD_XI12.XI19.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=1.125e-12 AS=9.375e-13
+ PD=3e-06 PS=2.75e-06
mXI12.XI20.MM27 N_XI12.XI20.NET31_XI12.XI20.MM27_d
+ N_XI12.XI20.NET35_XI12.XI20.MM27_g N_XI12.XI20.NET58_XI12.XI20.MM27_s
+ N_VDD_XI12.XI20.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=1.125e-12 AS=9.375e-13
+ PD=3e-06 PS=2.75e-06
mXI12.XI18.MM27 N_XI12.XI18.NET31_XI12.XI18.MM27_d
+ N_XI12.XI18.NET35_XI12.XI18.MM27_g N_XI12.XI18.NET58_XI12.XI18.MM27_s
+ N_VDD_XI12.XI18.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=1.125e-12 AS=9.375e-13
+ PD=3e-06 PS=2.75e-06
mXI12.XI17.MM27 N_XI12.XI17.NET31_XI12.XI17.MM27_d
+ N_XI12.XI17.NET35_XI12.XI17.MM27_g N_XI12.XI17.NET58_XI12.XI17.MM27_s
+ N_VDD_XI12.XI17.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=1.125e-12 AS=9.375e-13
+ PD=3e-06 PS=2.75e-06
mXI12.XI0.MM27 N_XI12.XI0.NET31_XI12.XI0.MM27_d N_XI12.XI0.NET35_XI12.XI0.MM27_g
+ N_XI12.XI0.NET58_XI12.XI0.MM27_s N_VDD_XI12.XI0.XI0.MM1_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.125e-12 AS=9.375e-13 PD=3e-06 PS=2.75e-06
mXI12.XI30.MM3 N_XI12.XI30.NET15_XI12.XI30.MM3_d
+ N_XI12.XI30.NET58_XI12.XI30.MM3_g N_VDD_XI12.XI30.MM3_s
+ N_VDD_XI12.XI30.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI12.XI29.MM3 N_XI12.XI29.NET15_XI12.XI29.MM3_d
+ N_XI12.XI29.NET58_XI12.XI29.MM3_g N_VDD_XI12.XI29.MM3_s
+ N_VDD_XI12.XI29.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI12.XI31.MM3 N_XI12.XI31.NET15_XI12.XI31.MM3_d
+ N_XI12.XI31.NET58_XI12.XI31.MM3_g N_VDD_XI12.XI31.MM3_s
+ N_VDD_XI12.XI31.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI12.XI28.MM3 N_XI12.XI28.NET15_XI12.XI28.MM3_d
+ N_XI12.XI28.NET58_XI12.XI28.MM3_g N_VDD_XI12.XI28.MM3_s
+ N_VDD_XI12.XI28.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI12.XI25.MM3 N_XI12.XI25.NET15_XI12.XI25.MM3_d
+ N_XI12.XI25.NET58_XI12.XI25.MM3_g N_VDD_XI12.XI25.MM3_s
+ N_VDD_XI12.XI25.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI12.XI26.MM3 N_XI12.XI26.NET15_XI12.XI26.MM3_d
+ N_XI12.XI26.NET58_XI12.XI26.MM3_g N_VDD_XI12.XI26.MM3_s
+ N_VDD_XI12.XI26.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI12.XI24.MM3 N_XI12.XI24.NET15_XI12.XI24.MM3_d
+ N_XI12.XI24.NET58_XI12.XI24.MM3_g N_VDD_XI12.XI24.MM3_s
+ N_VDD_XI12.XI24.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI12.XI27.MM3 N_XI12.XI27.NET15_XI12.XI27.MM3_d
+ N_XI12.XI27.NET58_XI12.XI27.MM3_g N_VDD_XI12.XI27.MM3_s
+ N_VDD_XI12.XI27.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI12.XI22.MM3 N_XI12.XI22.NET15_XI12.XI22.MM3_d
+ N_XI12.XI22.NET58_XI12.XI22.MM3_g N_VDD_XI12.XI22.MM3_s
+ N_VDD_XI12.XI22.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI12.XI21.MM3 N_XI12.XI21.NET15_XI12.XI21.MM3_d
+ N_XI12.XI21.NET58_XI12.XI21.MM3_g N_VDD_XI12.XI21.MM3_s
+ N_VDD_XI12.XI21.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI12.XI23.MM3 N_XI12.XI23.NET15_XI12.XI23.MM3_d
+ N_XI12.XI23.NET58_XI12.XI23.MM3_g N_VDD_XI12.XI23.MM3_s
+ N_VDD_XI12.XI23.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI12.XI19.MM3 N_XI12.XI19.NET15_XI12.XI19.MM3_d
+ N_XI12.XI19.NET58_XI12.XI19.MM3_g N_VDD_XI12.XI19.MM3_s
+ N_VDD_XI12.XI19.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI12.XI20.MM3 N_XI12.XI20.NET15_XI12.XI20.MM3_d
+ N_XI12.XI20.NET58_XI12.XI20.MM3_g N_VDD_XI12.XI20.MM3_s
+ N_VDD_XI12.XI20.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI12.XI18.MM3 N_XI12.XI18.NET15_XI12.XI18.MM3_d
+ N_XI12.XI18.NET58_XI12.XI18.MM3_g N_VDD_XI12.XI18.MM3_s
+ N_VDD_XI12.XI18.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI12.XI17.MM3 N_XI12.XI17.NET15_XI12.XI17.MM3_d
+ N_XI12.XI17.NET58_XI12.XI17.MM3_g N_VDD_XI12.XI17.MM3_s
+ N_VDD_XI12.XI17.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI12.XI0.MM3 N_XI12.XI0.NET15_XI12.XI0.MM3_d N_XI12.XI0.NET58_XI12.XI0.MM3_g
+ N_VDD_XI12.XI0.MM3_s N_VDD_XI12.XI0.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI12.XI30.MM1 N_XI12.XI30.NET54_XI12.XI30.MM1_d
+ N_XI12.XI30.NET15_XI12.XI30.MM1_g N_VDD_XI12.XI30.MM1_s
+ N_VDD_XI12.XI30.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI12.XI29.MM1 N_XI12.XI29.NET54_XI12.XI29.MM1_d
+ N_XI12.XI29.NET15_XI12.XI29.MM1_g N_VDD_XI12.XI29.MM1_s
+ N_VDD_XI12.XI29.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI12.XI31.MM1 N_XI12.XI31.NET54_XI12.XI31.MM1_d
+ N_XI12.XI31.NET15_XI12.XI31.MM1_g N_VDD_XI12.XI31.MM1_s
+ N_VDD_XI12.XI31.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI12.XI28.MM1 N_XI12.XI28.NET54_XI12.XI28.MM1_d
+ N_XI12.XI28.NET15_XI12.XI28.MM1_g N_VDD_XI12.XI28.MM1_s
+ N_VDD_XI12.XI28.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI12.XI25.MM1 N_XI12.XI25.NET54_XI12.XI25.MM1_d
+ N_XI12.XI25.NET15_XI12.XI25.MM1_g N_VDD_XI12.XI25.MM1_s
+ N_VDD_XI12.XI25.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI12.XI26.MM1 N_XI12.XI26.NET54_XI12.XI26.MM1_d
+ N_XI12.XI26.NET15_XI12.XI26.MM1_g N_VDD_XI12.XI26.MM1_s
+ N_VDD_XI12.XI26.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI12.XI24.MM1 N_XI12.XI24.NET54_XI12.XI24.MM1_d
+ N_XI12.XI24.NET15_XI12.XI24.MM1_g N_VDD_XI12.XI24.MM1_s
+ N_VDD_XI12.XI24.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI12.XI27.MM1 N_XI12.XI27.NET54_XI12.XI27.MM1_d
+ N_XI12.XI27.NET15_XI12.XI27.MM1_g N_VDD_XI12.XI27.MM1_s
+ N_VDD_XI12.XI27.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI12.XI22.MM1 N_XI12.XI22.NET54_XI12.XI22.MM1_d
+ N_XI12.XI22.NET15_XI12.XI22.MM1_g N_VDD_XI12.XI22.MM1_s
+ N_VDD_XI12.XI22.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI12.XI21.MM1 N_XI12.XI21.NET54_XI12.XI21.MM1_d
+ N_XI12.XI21.NET15_XI12.XI21.MM1_g N_VDD_XI12.XI21.MM1_s
+ N_VDD_XI12.XI21.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI12.XI23.MM1 N_XI12.XI23.NET54_XI12.XI23.MM1_d
+ N_XI12.XI23.NET15_XI12.XI23.MM1_g N_VDD_XI12.XI23.MM1_s
+ N_VDD_XI12.XI23.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI12.XI19.MM1 N_XI12.XI19.NET54_XI12.XI19.MM1_d
+ N_XI12.XI19.NET15_XI12.XI19.MM1_g N_VDD_XI12.XI19.MM1_s
+ N_VDD_XI12.XI19.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI12.XI20.MM1 N_XI12.XI20.NET54_XI12.XI20.MM1_d
+ N_XI12.XI20.NET15_XI12.XI20.MM1_g N_VDD_XI12.XI20.MM1_s
+ N_VDD_XI12.XI20.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI12.XI18.MM1 N_XI12.XI18.NET54_XI12.XI18.MM1_d
+ N_XI12.XI18.NET15_XI12.XI18.MM1_g N_VDD_XI12.XI18.MM1_s
+ N_VDD_XI12.XI18.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI12.XI17.MM1 N_XI12.XI17.NET54_XI12.XI17.MM1_d
+ N_XI12.XI17.NET15_XI12.XI17.MM1_g N_VDD_XI12.XI17.MM1_s
+ N_VDD_XI12.XI17.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI12.XI0.MM1 N_XI12.XI0.NET54_XI12.XI0.MM1_d N_XI12.XI0.NET15_XI12.XI0.MM1_g
+ N_VDD_XI12.XI0.MM1_s N_VDD_XI12.XI0.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI12.XI30.MM35 N_XI12.XI30.NET58_XI12.XI30.MM35_d
+ N_XI12.XI30.CLKB_XI12.XI30.MM35_g N_XI12.XI30.NET54_XI12.XI30.MM35_s
+ N_VDD_XI12.XI30.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI12.XI29.MM35 N_XI12.XI29.NET58_XI12.XI29.MM35_d
+ N_XI12.XI29.CLKB_XI12.XI29.MM35_g N_XI12.XI29.NET54_XI12.XI29.MM35_s
+ N_VDD_XI12.XI29.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI12.XI31.MM35 N_XI12.XI31.NET58_XI12.XI31.MM35_d
+ N_XI12.XI31.CLKB_XI12.XI31.MM35_g N_XI12.XI31.NET54_XI12.XI31.MM35_s
+ N_VDD_XI12.XI31.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI12.XI28.MM35 N_XI12.XI28.NET58_XI12.XI28.MM35_d
+ N_XI12.XI28.CLKB_XI12.XI28.MM35_g N_XI12.XI28.NET54_XI12.XI28.MM35_s
+ N_VDD_XI12.XI28.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI12.XI25.MM35 N_XI12.XI25.NET58_XI12.XI25.MM35_d
+ N_XI12.XI25.CLKB_XI12.XI25.MM35_g N_XI12.XI25.NET54_XI12.XI25.MM35_s
+ N_VDD_XI12.XI25.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI12.XI26.MM35 N_XI12.XI26.NET58_XI12.XI26.MM35_d
+ N_XI12.XI26.CLKB_XI12.XI26.MM35_g N_XI12.XI26.NET54_XI12.XI26.MM35_s
+ N_VDD_XI12.XI26.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI12.XI24.MM35 N_XI12.XI24.NET58_XI12.XI24.MM35_d
+ N_XI12.XI24.CLKB_XI12.XI24.MM35_g N_XI12.XI24.NET54_XI12.XI24.MM35_s
+ N_VDD_XI12.XI24.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI12.XI27.MM35 N_XI12.XI27.NET58_XI12.XI27.MM35_d
+ N_XI12.XI27.CLKB_XI12.XI27.MM35_g N_XI12.XI27.NET54_XI12.XI27.MM35_s
+ N_VDD_XI12.XI27.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI12.XI22.MM35 N_XI12.XI22.NET58_XI12.XI22.MM35_d
+ N_XI12.XI22.CLKB_XI12.XI22.MM35_g N_XI12.XI22.NET54_XI12.XI22.MM35_s
+ N_VDD_XI12.XI22.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI12.XI21.MM35 N_XI12.XI21.NET58_XI12.XI21.MM35_d
+ N_XI12.XI21.CLKB_XI12.XI21.MM35_g N_XI12.XI21.NET54_XI12.XI21.MM35_s
+ N_VDD_XI12.XI21.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI12.XI23.MM35 N_XI12.XI23.NET58_XI12.XI23.MM35_d
+ N_XI12.XI23.CLKB_XI12.XI23.MM35_g N_XI12.XI23.NET54_XI12.XI23.MM35_s
+ N_VDD_XI12.XI23.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI12.XI19.MM35 N_XI12.XI19.NET58_XI12.XI19.MM35_d
+ N_XI12.XI19.CLKB_XI12.XI19.MM35_g N_XI12.XI19.NET54_XI12.XI19.MM35_s
+ N_VDD_XI12.XI19.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI12.XI20.MM35 N_XI12.XI20.NET58_XI12.XI20.MM35_d
+ N_XI12.XI20.CLKB_XI12.XI20.MM35_g N_XI12.XI20.NET54_XI12.XI20.MM35_s
+ N_VDD_XI12.XI20.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI12.XI18.MM35 N_XI12.XI18.NET58_XI12.XI18.MM35_d
+ N_XI12.XI18.CLKB_XI12.XI18.MM35_g N_XI12.XI18.NET54_XI12.XI18.MM35_s
+ N_VDD_XI12.XI18.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI12.XI17.MM35 N_XI12.XI17.NET58_XI12.XI17.MM35_d
+ N_XI12.XI17.CLKB_XI12.XI17.MM35_g N_XI12.XI17.NET54_XI12.XI17.MM35_s
+ N_VDD_XI12.XI17.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI12.XI0.MM35 N_XI12.XI0.NET58_XI12.XI0.MM35_d N_XI12.XI0.CLKB_XI12.XI0.MM35_g
+ N_XI12.XI0.NET54_XI12.XI0.MM35_s N_VDD_XI12.XI0.XI0.MM1_b P_18 L=1.8e-07
+ W=1.5e-06 AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI12.XI30.MM37 N_XI12.XI30.NET15_XI12.XI30.MM37_d
+ N_XI12.XI30.CLKB_XI12.XI30.MM37_g N_XI12.XI30.NET14_XI12.XI30.MM37_s
+ N_VDD_XI12.XI30.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=1.125e-12 AS=9.375e-13
+ PD=3e-06 PS=2.75e-06
mXI12.XI29.MM37 N_XI12.XI29.NET15_XI12.XI29.MM37_d
+ N_XI12.XI29.CLKB_XI12.XI29.MM37_g N_XI12.XI29.NET14_XI12.XI29.MM37_s
+ N_VDD_XI12.XI29.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=1.125e-12 AS=9.375e-13
+ PD=3e-06 PS=2.75e-06
mXI12.XI31.MM37 N_XI12.XI31.NET15_XI12.XI31.MM37_d
+ N_XI12.XI31.CLKB_XI12.XI31.MM37_g N_XI12.XI31.NET14_XI12.XI31.MM37_s
+ N_VDD_XI12.XI31.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=1.125e-12 AS=9.375e-13
+ PD=3e-06 PS=2.75e-06
mXI12.XI28.MM37 N_XI12.XI28.NET15_XI12.XI28.MM37_d
+ N_XI12.XI28.CLKB_XI12.XI28.MM37_g N_XI12.XI28.NET14_XI12.XI28.MM37_s
+ N_VDD_XI12.XI28.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=1.125e-12 AS=9.375e-13
+ PD=3e-06 PS=2.75e-06
mXI12.XI25.MM37 N_XI12.XI25.NET15_XI12.XI25.MM37_d
+ N_XI12.XI25.CLKB_XI12.XI25.MM37_g N_XI12.XI25.NET14_XI12.XI25.MM37_s
+ N_VDD_XI12.XI25.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=1.125e-12 AS=9.375e-13
+ PD=3e-06 PS=2.75e-06
mXI12.XI26.MM37 N_XI12.XI26.NET15_XI12.XI26.MM37_d
+ N_XI12.XI26.CLKB_XI12.XI26.MM37_g N_XI12.XI26.NET14_XI12.XI26.MM37_s
+ N_VDD_XI12.XI26.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=1.125e-12 AS=9.375e-13
+ PD=3e-06 PS=2.75e-06
mXI12.XI24.MM37 N_XI12.XI24.NET15_XI12.XI24.MM37_d
+ N_XI12.XI24.CLKB_XI12.XI24.MM37_g N_XI12.XI24.NET14_XI12.XI24.MM37_s
+ N_VDD_XI12.XI24.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=1.125e-12 AS=9.375e-13
+ PD=3e-06 PS=2.75e-06
mXI12.XI27.MM37 N_XI12.XI27.NET15_XI12.XI27.MM37_d
+ N_XI12.XI27.CLKB_XI12.XI27.MM37_g N_XI12.XI27.NET14_XI12.XI27.MM37_s
+ N_VDD_XI12.XI27.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=1.125e-12 AS=9.375e-13
+ PD=3e-06 PS=2.75e-06
mXI12.XI22.MM37 N_XI12.XI22.NET15_XI12.XI22.MM37_d
+ N_XI12.XI22.CLKB_XI12.XI22.MM37_g N_XI12.XI22.NET14_XI12.XI22.MM37_s
+ N_VDD_XI12.XI22.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=1.125e-12 AS=9.375e-13
+ PD=3e-06 PS=2.75e-06
mXI12.XI21.MM37 N_XI12.XI21.NET15_XI12.XI21.MM37_d
+ N_XI12.XI21.CLKB_XI12.XI21.MM37_g N_XI12.XI21.NET14_XI12.XI21.MM37_s
+ N_VDD_XI12.XI21.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=1.125e-12 AS=9.375e-13
+ PD=3e-06 PS=2.75e-06
mXI12.XI23.MM37 N_XI12.XI23.NET15_XI12.XI23.MM37_d
+ N_XI12.XI23.CLKB_XI12.XI23.MM37_g N_XI12.XI23.NET14_XI12.XI23.MM37_s
+ N_VDD_XI12.XI23.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=1.125e-12 AS=9.375e-13
+ PD=3e-06 PS=2.75e-06
mXI12.XI19.MM37 N_XI12.XI19.NET15_XI12.XI19.MM37_d
+ N_XI12.XI19.CLKB_XI12.XI19.MM37_g N_XI12.XI19.NET14_XI12.XI19.MM37_s
+ N_VDD_XI12.XI19.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=1.125e-12 AS=9.375e-13
+ PD=3e-06 PS=2.75e-06
mXI12.XI20.MM37 N_XI12.XI20.NET15_XI12.XI20.MM37_d
+ N_XI12.XI20.CLKB_XI12.XI20.MM37_g N_XI12.XI20.NET14_XI12.XI20.MM37_s
+ N_VDD_XI12.XI20.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=1.125e-12 AS=9.375e-13
+ PD=3e-06 PS=2.75e-06
mXI12.XI18.MM37 N_XI12.XI18.NET15_XI12.XI18.MM37_d
+ N_XI12.XI18.CLKB_XI12.XI18.MM37_g N_XI12.XI18.NET14_XI12.XI18.MM37_s
+ N_VDD_XI12.XI18.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=1.125e-12 AS=9.375e-13
+ PD=3e-06 PS=2.75e-06
mXI12.XI17.MM37 N_XI12.XI17.NET15_XI12.XI17.MM37_d
+ N_XI12.XI17.CLKB_XI12.XI17.MM37_g N_XI12.XI17.NET14_XI12.XI17.MM37_s
+ N_VDD_XI12.XI17.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=1.125e-12 AS=9.375e-13
+ PD=3e-06 PS=2.75e-06
mXI12.XI0.MM37 N_XI12.XI0.NET15_XI12.XI0.MM37_d N_XI12.XI0.CLKB_XI12.XI0.MM37_g
+ N_XI12.XI0.NET14_XI12.XI0.MM37_s N_VDD_XI12.XI0.XI0.MM1_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.125e-12 AS=9.375e-13 PD=3e-06 PS=2.75e-06
mXI12.XI30.MM13 N_MIN15_XI12.XI30.MM13_d N_XI12.XI30.NET14_XI12.XI30.MM13_g
+ N_VDD_XI12.XI30.MM13_s N_VDD_XI12.XI30.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI12.XI29.MM13 N_MIN14_XI12.XI29.MM13_d N_XI12.XI29.NET14_XI12.XI29.MM13_g
+ N_VDD_XI12.XI29.MM13_s N_VDD_XI12.XI29.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI12.XI31.MM13 N_MIN13_XI12.XI31.MM13_d N_XI12.XI31.NET14_XI12.XI31.MM13_g
+ N_VDD_XI12.XI31.MM13_s N_VDD_XI12.XI31.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI12.XI28.MM13 N_MIN12_XI12.XI28.MM13_d N_XI12.XI28.NET14_XI12.XI28.MM13_g
+ N_VDD_XI12.XI28.MM13_s N_VDD_XI12.XI28.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI12.XI25.MM13 N_MIN11_XI12.XI25.MM13_d N_XI12.XI25.NET14_XI12.XI25.MM13_g
+ N_VDD_XI12.XI25.MM13_s N_VDD_XI12.XI25.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI12.XI26.MM13 N_MIN10_XI12.XI26.MM13_d N_XI12.XI26.NET14_XI12.XI26.MM13_g
+ N_VDD_XI12.XI26.MM13_s N_VDD_XI12.XI26.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI12.XI24.MM13 N_MIN9_XI12.XI24.MM13_d N_XI12.XI24.NET14_XI12.XI24.MM13_g
+ N_VDD_XI12.XI24.MM13_s N_VDD_XI12.XI24.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI12.XI27.MM13 N_MIN8_XI12.XI27.MM13_d N_XI12.XI27.NET14_XI12.XI27.MM13_g
+ N_VDD_XI12.XI27.MM13_s N_VDD_XI12.XI27.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI12.XI22.MM13 N_MIN7_XI12.XI22.MM13_d N_XI12.XI22.NET14_XI12.XI22.MM13_g
+ N_VDD_XI12.XI22.MM13_s N_VDD_XI12.XI22.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI12.XI21.MM13 N_MIN6_XI12.XI21.MM13_d N_XI12.XI21.NET14_XI12.XI21.MM13_g
+ N_VDD_XI12.XI21.MM13_s N_VDD_XI12.XI21.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI12.XI23.MM13 N_MIN5_XI12.XI23.MM13_d N_XI12.XI23.NET14_XI12.XI23.MM13_g
+ N_VDD_XI12.XI23.MM13_s N_VDD_XI12.XI23.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI12.XI19.MM13 N_MIN4_XI12.XI19.MM13_d N_XI12.XI19.NET14_XI12.XI19.MM13_g
+ N_VDD_XI12.XI19.MM13_s N_VDD_XI12.XI19.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI12.XI20.MM13 N_MIN3_XI12.XI20.MM13_d N_XI12.XI20.NET14_XI12.XI20.MM13_g
+ N_VDD_XI12.XI20.MM13_s N_VDD_XI12.XI20.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI12.XI18.MM13 N_MIN2_XI12.XI18.MM13_d N_XI12.XI18.NET14_XI12.XI18.MM13_g
+ N_VDD_XI12.XI18.MM13_s N_VDD_XI12.XI18.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI12.XI17.MM13 N_MIN1_XI12.XI17.MM13_d N_XI12.XI17.NET14_XI12.XI17.MM13_g
+ N_VDD_XI12.XI17.MM13_s N_VDD_XI12.XI17.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI12.XI0.MM13 N_MIN0_XI12.XI0.MM13_d N_XI12.XI0.NET14_XI12.XI0.MM13_g
+ N_VDD_XI12.XI0.MM13_s N_VDD_XI12.XI0.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI12.XI30.MM14 N_XI12.BAR_Q16_XI12.XI30.MM14_d N_MIN15_XI12.XI30.MM14_g
+ N_VDD_XI12.XI30.MM14_s N_VDD_XI12.XI30.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI12.XI29.MM14 N_XI12.BAR_Q15_XI12.XI29.MM14_d N_MIN14_XI12.XI29.MM14_g
+ N_VDD_XI12.XI29.MM14_s N_VDD_XI12.XI29.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI12.XI31.MM14 N_XI12.BAR_Q14_XI12.XI31.MM14_d N_MIN13_XI12.XI31.MM14_g
+ N_VDD_XI12.XI31.MM14_s N_VDD_XI12.XI31.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI12.XI28.MM14 N_XI12.BAR_Q13_XI12.XI28.MM14_d N_MIN12_XI12.XI28.MM14_g
+ N_VDD_XI12.XI28.MM14_s N_VDD_XI12.XI28.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI12.XI25.MM14 N_XI12.BAR_Q12_XI12.XI25.MM14_d N_MIN11_XI12.XI25.MM14_g
+ N_VDD_XI12.XI25.MM14_s N_VDD_XI12.XI25.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI12.XI26.MM14 N_XI12.BAR_Q11_XI12.XI26.MM14_d N_MIN10_XI12.XI26.MM14_g
+ N_VDD_XI12.XI26.MM14_s N_VDD_XI12.XI26.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI12.XI24.MM14 N_XI12.BAR_Q10_XI12.XI24.MM14_d N_MIN9_XI12.XI24.MM14_g
+ N_VDD_XI12.XI24.MM14_s N_VDD_XI12.XI24.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI12.XI27.MM14 N_XI12.BAR_Q9_XI12.XI27.MM14_d N_MIN8_XI12.XI27.MM14_g
+ N_VDD_XI12.XI27.MM14_s N_VDD_XI12.XI27.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI12.XI22.MM14 N_XI12.BAR_Q8_XI12.XI22.MM14_d N_MIN7_XI12.XI22.MM14_g
+ N_VDD_XI12.XI22.MM14_s N_VDD_XI12.XI22.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI12.XI21.MM14 N_XI12.BAR_Q7_XI12.XI21.MM14_d N_MIN6_XI12.XI21.MM14_g
+ N_VDD_XI12.XI21.MM14_s N_VDD_XI12.XI21.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI12.XI23.MM14 N_XI12.BAR_Q6_XI12.XI23.MM14_d N_MIN5_XI12.XI23.MM14_g
+ N_VDD_XI12.XI23.MM14_s N_VDD_XI12.XI23.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI12.XI19.MM14 N_XI12.BAR_Q5_XI12.XI19.MM14_d N_MIN4_XI12.XI19.MM14_g
+ N_VDD_XI12.XI19.MM14_s N_VDD_XI12.XI19.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI12.XI20.MM14 N_XI12.BAR_Q4_XI12.XI20.MM14_d N_MIN3_XI12.XI20.MM14_g
+ N_VDD_XI12.XI20.MM14_s N_VDD_XI12.XI20.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI12.XI18.MM14 N_XI12.BAR_Q3_XI12.XI18.MM14_d N_MIN2_XI12.XI18.MM14_g
+ N_VDD_XI12.XI18.MM14_s N_VDD_XI12.XI18.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI12.XI17.MM14 N_XI12.BAR_Q2_XI12.XI17.MM14_d N_MIN1_XI12.XI17.MM14_g
+ N_VDD_XI12.XI17.MM14_s N_VDD_XI12.XI17.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI12.XI0.MM14 N_XI12.BAR_Q1_XI12.XI0.MM14_d N_MIN0_XI12.XI0.MM14_g
+ N_VDD_XI12.XI0.MM14_s N_VDD_XI12.XI0.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI12.XI30.MM39 N_XI12.XI30.NET14_XI12.XI30.MM39_d
+ N_XI12.XI30.NET35_XI12.XI30.MM39_g N_XI12.BAR_Q16_XI12.XI30.MM39_s
+ N_VDD_XI12.XI30.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI12.XI29.MM39 N_XI12.XI29.NET14_XI12.XI29.MM39_d
+ N_XI12.XI29.NET35_XI12.XI29.MM39_g N_XI12.BAR_Q15_XI12.XI29.MM39_s
+ N_VDD_XI12.XI29.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI12.XI31.MM39 N_XI12.XI31.NET14_XI12.XI31.MM39_d
+ N_XI12.XI31.NET35_XI12.XI31.MM39_g N_XI12.BAR_Q14_XI12.XI31.MM39_s
+ N_VDD_XI12.XI31.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI12.XI28.MM39 N_XI12.XI28.NET14_XI12.XI28.MM39_d
+ N_XI12.XI28.NET35_XI12.XI28.MM39_g N_XI12.BAR_Q13_XI12.XI28.MM39_s
+ N_VDD_XI12.XI28.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI12.XI25.MM39 N_XI12.XI25.NET14_XI12.XI25.MM39_d
+ N_XI12.XI25.NET35_XI12.XI25.MM39_g N_XI12.BAR_Q12_XI12.XI25.MM39_s
+ N_VDD_XI12.XI25.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI12.XI26.MM39 N_XI12.XI26.NET14_XI12.XI26.MM39_d
+ N_XI12.XI26.NET35_XI12.XI26.MM39_g N_XI12.BAR_Q11_XI12.XI26.MM39_s
+ N_VDD_XI12.XI26.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI12.XI24.MM39 N_XI12.XI24.NET14_XI12.XI24.MM39_d
+ N_XI12.XI24.NET35_XI12.XI24.MM39_g N_XI12.BAR_Q10_XI12.XI24.MM39_s
+ N_VDD_XI12.XI24.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI12.XI27.MM39 N_XI12.XI27.NET14_XI12.XI27.MM39_d
+ N_XI12.XI27.NET35_XI12.XI27.MM39_g N_XI12.BAR_Q9_XI12.XI27.MM39_s
+ N_VDD_XI12.XI27.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI12.XI22.MM39 N_XI12.XI22.NET14_XI12.XI22.MM39_d
+ N_XI12.XI22.NET35_XI12.XI22.MM39_g N_XI12.BAR_Q8_XI12.XI22.MM39_s
+ N_VDD_XI12.XI22.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI12.XI21.MM39 N_XI12.XI21.NET14_XI12.XI21.MM39_d
+ N_XI12.XI21.NET35_XI12.XI21.MM39_g N_XI12.BAR_Q7_XI12.XI21.MM39_s
+ N_VDD_XI12.XI21.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI12.XI23.MM39 N_XI12.XI23.NET14_XI12.XI23.MM39_d
+ N_XI12.XI23.NET35_XI12.XI23.MM39_g N_XI12.BAR_Q6_XI12.XI23.MM39_s
+ N_VDD_XI12.XI23.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI12.XI19.MM39 N_XI12.XI19.NET14_XI12.XI19.MM39_d
+ N_XI12.XI19.NET35_XI12.XI19.MM39_g N_XI12.BAR_Q5_XI12.XI19.MM39_s
+ N_VDD_XI12.XI19.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI12.XI20.MM39 N_XI12.XI20.NET14_XI12.XI20.MM39_d
+ N_XI12.XI20.NET35_XI12.XI20.MM39_g N_XI12.BAR_Q4_XI12.XI20.MM39_s
+ N_VDD_XI12.XI20.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI12.XI18.MM39 N_XI12.XI18.NET14_XI12.XI18.MM39_d
+ N_XI12.XI18.NET35_XI12.XI18.MM39_g N_XI12.BAR_Q3_XI12.XI18.MM39_s
+ N_VDD_XI12.XI18.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI12.XI17.MM39 N_XI12.XI17.NET14_XI12.XI17.MM39_d
+ N_XI12.XI17.NET35_XI12.XI17.MM39_g N_XI12.BAR_Q2_XI12.XI17.MM39_s
+ N_VDD_XI12.XI17.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI12.XI0.MM39 N_XI12.XI0.NET14_XI12.XI0.MM39_d N_XI12.XI0.NET35_XI12.XI0.MM39_g
+ N_XI12.BAR_Q1_XI12.XI0.MM39_s N_VDD_XI12.XI0.XI0.MM1_b P_18 L=1.8e-07
+ W=1.5e-06 AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI1.XI134.XI9.MM1 N_XI1.XI134.NET43_XI1.XI134.XI9.MM1_d
+ N_NET628_XI1.XI134.XI9.MM1_g N_VDD_XI1.XI134.XI9.MM1_s
+ N_VDD_XI1.XI134.XI9.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI1.XI153.XI1.MM3 N_XI1.XI153.NET6_XI1.XI153.XI1.MM3_d
+ N_NET629_XI1.XI153.XI1.MM3_g N_VDD_XI1.XI153.XI1.MM3_s
+ N_VDD_XI1.XI153.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.35e-13
+ PD=7.4e-07 PS=2.48e-06
mXI1.XI154.XI1.MM3 N_XI1.XI154.NET6_XI1.XI154.XI1.MM3_d
+ N_NET630_XI1.XI154.XI1.MM3_g N_VDD_XI1.XI154.XI1.MM3_s
+ N_VDD_XI1.XI154.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.35e-13
+ PD=7.4e-07 PS=2.48e-06
mXI1.XI157.XI1.MM3 N_XI1.XI157.NET6_XI1.XI157.XI1.MM3_d
+ N_NET631_XI1.XI157.XI1.MM3_g N_VDD_XI1.XI157.XI1.MM3_s
+ N_VDD_XI1.XI157.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.35e-13
+ PD=7.4e-07 PS=2.48e-06
mXI1.XI156.XI1.MM3 N_XI1.XI156.NET6_XI1.XI156.XI1.MM3_d
+ N_NET632_XI1.XI156.XI1.MM3_g N_VDD_XI1.XI156.XI1.MM3_s
+ N_VDD_XI1.XI156.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.35e-13
+ PD=7.4e-07 PS=2.48e-06
mXI1.XI155.XI1.MM3 N_XI1.XI155.NET6_XI1.XI155.XI1.MM3_d
+ N_NET633_XI1.XI155.XI1.MM3_g N_VDD_XI1.XI155.XI1.MM3_s
+ N_VDD_XI1.XI155.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.35e-13
+ PD=7.4e-07 PS=2.48e-06
mXI1.XI133.XI1.MM3 N_XI1.XI133.NET6_XI1.XI133.XI1.MM3_d
+ N_NET634_XI1.XI133.XI1.MM3_g N_VDD_XI1.XI133.XI1.MM3_s
+ N_VDD_XI1.XI133.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.35e-13
+ PD=7.4e-07 PS=2.48e-06
mXI1.XI132.XI1.MM3 N_XI1.XI132.NET6_XI1.XI132.XI1.MM3_d
+ N_NET635_XI1.XI132.XI1.MM3_g N_VDD_XI1.XI132.XI1.MM3_s
+ N_VDD_XI1.XI132.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.35e-13
+ PD=7.4e-07 PS=2.48e-06
mXI1.XI131.XI1.MM3 N_XI1.XI131.NET6_XI1.XI131.XI1.MM3_d
+ N_NET636_XI1.XI131.XI1.MM3_g N_VDD_XI1.XI131.XI1.MM3_s
+ N_VDD_XI1.XI131.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.35e-13
+ PD=7.4e-07 PS=2.48e-06
mXI1.XI111.XI1.MM3 N_XI1.XI111.NET6_XI1.XI111.XI1.MM3_d
+ N_NET637_XI1.XI111.XI1.MM3_g N_VDD_XI1.XI111.XI1.MM3_s
+ N_VDD_XI1.XI111.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.35e-13
+ PD=7.4e-07 PS=2.48e-06
mXI1.XI110.XI1.MM3 N_XI1.XI110.NET6_XI1.XI110.XI1.MM3_d
+ N_NET638_XI1.XI110.XI1.MM3_g N_VDD_XI1.XI110.XI1.MM3_s
+ N_VDD_XI1.XI110.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.35e-13
+ PD=7.4e-07 PS=2.48e-06
mXI1.XI103.XI1.MM3 N_XI1.XI103.NET6_XI1.XI103.XI1.MM3_d
+ N_NET639_XI1.XI103.XI1.MM3_g N_VDD_XI1.XI103.XI1.MM3_s
+ N_VDD_XI1.XI103.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.35e-13
+ PD=7.4e-07 PS=2.48e-06
mXI1.XI102.XI1.MM3 N_XI1.XI102.NET6_XI1.XI102.XI1.MM3_d
+ N_NET640_XI1.XI102.XI1.MM3_g N_VDD_XI1.XI102.XI1.MM3_s
+ N_VDD_XI1.XI102.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.35e-13
+ PD=7.4e-07 PS=2.48e-06
mXI1.XI88.XI1.MM3 N_XI1.XI88.NET6_XI1.XI88.XI1.MM3_d N_NET641_XI1.XI88.XI1.MM3_g
+ N_VDD_XI1.XI88.XI1.MM3_s N_VDD_XI1.XI88.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=5.55e-13 AS=7.35e-13 PD=7.4e-07 PS=2.48e-06
mXI1.XI82.XI1.MM3 N_XI1.XI82.NET6_XI1.XI82.XI1.MM3_d N_NET642_XI1.XI82.XI1.MM3_g
+ N_VDD_XI1.XI82.XI1.MM3_s N_VDD_XI1.XI82.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=5.55e-13 AS=7.35e-13 PD=7.4e-07 PS=2.48e-06
mXI1.XI10.XI1.MM3 N_XI1.XI10.NET6_XI1.XI10.XI1.MM3_d N_NET643_XI1.XI10.XI1.MM3_g
+ N_VDD_XI1.XI10.XI1.MM3_s N_VDD_XI1.XI10.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=5.55e-13 AS=7.35e-13 PD=7.4e-07 PS=2.48e-06
mXI3.MM1 N_NET01249_XI3.MM1_d N_NET0855_XI3.MM1_g N_VDD_XI3.MM1_s
+ N_VDD_XI3.MM1_b P_18 L=1.8e-07 W=9e-06 AD=4.41e-12 AS=4.41e-12 PD=9.98e-06
+ PS=9.98e-06
mXI1.XI153.XI1.MM1 N_XI1.XI153.NET6_XI1.XI153.XI1.MM1_d
+ N_MAX14_XI1.XI153.XI1.MM1_g N_VDD_XI1.XI153.XI1.MM1_s
+ N_VDD_XI1.XI153.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.65e-13
+ PD=7.4e-07 PS=2.52e-06
mXI1.XI154.XI1.MM1 N_XI1.XI154.NET6_XI1.XI154.XI1.MM1_d
+ N_MAX13_XI1.XI154.XI1.MM1_g N_VDD_XI1.XI154.XI1.MM1_s
+ N_VDD_XI1.XI154.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.65e-13
+ PD=7.4e-07 PS=2.52e-06
mXI1.XI157.XI1.MM1 N_XI1.XI157.NET6_XI1.XI157.XI1.MM1_d
+ N_MAX12_XI1.XI157.XI1.MM1_g N_VDD_XI1.XI157.XI1.MM1_s
+ N_VDD_XI1.XI157.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.65e-13
+ PD=7.4e-07 PS=2.52e-06
mXI1.XI156.XI1.MM1 N_XI1.XI156.NET6_XI1.XI156.XI1.MM1_d
+ N_MAX11_XI1.XI156.XI1.MM1_g N_VDD_XI1.XI156.XI1.MM1_s
+ N_VDD_XI1.XI156.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.65e-13
+ PD=7.4e-07 PS=2.52e-06
mXI1.XI155.XI1.MM1 N_XI1.XI155.NET6_XI1.XI155.XI1.MM1_d
+ N_MAX10_XI1.XI155.XI1.MM1_g N_VDD_XI1.XI155.XI1.MM1_s
+ N_VDD_XI1.XI155.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.65e-13
+ PD=7.4e-07 PS=2.52e-06
mXI1.XI133.XI1.MM1 N_XI1.XI133.NET6_XI1.XI133.XI1.MM1_d
+ N_MAX9_XI1.XI133.XI1.MM1_g N_VDD_XI1.XI133.XI1.MM1_s N_VDD_XI1.XI133.XI1.MM3_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.65e-13 PD=7.4e-07 PS=2.52e-06
mXI1.XI132.XI1.MM1 N_XI1.XI132.NET6_XI1.XI132.XI1.MM1_d
+ N_MAX8_XI1.XI132.XI1.MM1_g N_VDD_XI1.XI132.XI1.MM1_s N_VDD_XI1.XI132.XI1.MM3_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.65e-13 PD=7.4e-07 PS=2.52e-06
mXI1.XI131.XI1.MM1 N_XI1.XI131.NET6_XI1.XI131.XI1.MM1_d
+ N_MAX7_XI1.XI131.XI1.MM1_g N_VDD_XI1.XI131.XI1.MM1_s N_VDD_XI1.XI131.XI1.MM3_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.65e-13 PD=7.4e-07 PS=2.52e-06
mXI1.XI111.XI1.MM1 N_XI1.XI111.NET6_XI1.XI111.XI1.MM1_d
+ N_MAX6_XI1.XI111.XI1.MM1_g N_VDD_XI1.XI111.XI1.MM1_s N_VDD_XI1.XI111.XI1.MM3_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.65e-13 PD=7.4e-07 PS=2.52e-06
mXI1.XI110.XI1.MM1 N_XI1.XI110.NET6_XI1.XI110.XI1.MM1_d
+ N_MAX5_XI1.XI110.XI1.MM1_g N_VDD_XI1.XI110.XI1.MM1_s N_VDD_XI1.XI110.XI1.MM3_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.65e-13 PD=7.4e-07 PS=2.52e-06
mXI1.XI103.XI1.MM1 N_XI1.XI103.NET6_XI1.XI103.XI1.MM1_d
+ N_MAX4_XI1.XI103.XI1.MM1_g N_VDD_XI1.XI103.XI1.MM1_s N_VDD_XI1.XI103.XI1.MM3_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.65e-13 PD=7.4e-07 PS=2.52e-06
mXI1.XI102.XI1.MM1 N_XI1.XI102.NET6_XI1.XI102.XI1.MM1_d
+ N_MAX3_XI1.XI102.XI1.MM1_g N_VDD_XI1.XI102.XI1.MM1_s N_VDD_XI1.XI102.XI1.MM3_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.65e-13 PD=7.4e-07 PS=2.52e-06
mXI1.XI88.XI1.MM1 N_XI1.XI88.NET6_XI1.XI88.XI1.MM1_d N_MAX2_XI1.XI88.XI1.MM1_g
+ N_VDD_XI1.XI88.XI1.MM1_s N_VDD_XI1.XI88.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=5.55e-13 AS=7.65e-13 PD=7.4e-07 PS=2.52e-06
mXI1.XI82.XI1.MM1 N_XI1.XI82.NET6_XI1.XI82.XI1.MM1_d N_MAX1_XI1.XI82.XI1.MM1_g
+ N_VDD_XI1.XI82.XI1.MM1_s N_VDD_XI1.XI82.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=5.55e-13 AS=7.65e-13 PD=7.4e-07 PS=2.52e-06
mXI1.XI10.XI1.MM1 N_XI1.XI10.NET6_XI1.XI10.XI1.MM1_d N_MAX0_XI1.XI10.XI1.MM1_g
+ N_VDD_XI1.XI10.XI1.MM1_s N_VDD_XI1.XI10.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=5.55e-13 AS=7.65e-13 PD=7.4e-07 PS=2.52e-06
mXI1.XI134.MM5 N_XI1.XI134.NET25_XI1.XI134.MM5_d
+ N_XI1.XI134.NET43_XI1.XI134.MM5_g N_VDD_XI1.XI134.MM5_s
+ N_VDD_XI1.XI134.XI9.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=6.7125e-13 AS=9.675e-13
+ PD=8.95e-07 PS=2.79e-06
mXI1.XI153.XI0.MM1 N_XI1.G15_XI1.XI153.XI0.MM1_d
+ N_XI1.XI153.NET6_XI1.XI153.XI0.MM1_g N_VDD_XI1.XI153.XI0.MM1_s
+ N_VDD_XI1.XI153.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI1.XI154.XI0.MM1 N_XI1.G14_XI1.XI154.XI0.MM1_d
+ N_XI1.XI154.NET6_XI1.XI154.XI0.MM1_g N_VDD_XI1.XI154.XI0.MM1_s
+ N_VDD_XI1.XI154.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI1.XI157.XI0.MM1 N_XI1.G13_XI1.XI157.XI0.MM1_d
+ N_XI1.XI157.NET6_XI1.XI157.XI0.MM1_g N_VDD_XI1.XI157.XI0.MM1_s
+ N_VDD_XI1.XI157.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI1.XI156.XI0.MM1 N_XI1.G12_XI1.XI156.XI0.MM1_d
+ N_XI1.XI156.NET6_XI1.XI156.XI0.MM1_g N_VDD_XI1.XI156.XI0.MM1_s
+ N_VDD_XI1.XI156.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI1.XI155.XI0.MM1 N_XI1.G11_XI1.XI155.XI0.MM1_d
+ N_XI1.XI155.NET6_XI1.XI155.XI0.MM1_g N_VDD_XI1.XI155.XI0.MM1_s
+ N_VDD_XI1.XI155.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI1.XI133.XI0.MM1 N_XI1.G10_XI1.XI133.XI0.MM1_d
+ N_XI1.XI133.NET6_XI1.XI133.XI0.MM1_g N_VDD_XI1.XI133.XI0.MM1_s
+ N_VDD_XI1.XI133.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI1.XI132.XI0.MM1 N_XI1.G9_XI1.XI132.XI0.MM1_d
+ N_XI1.XI132.NET6_XI1.XI132.XI0.MM1_g N_VDD_XI1.XI132.XI0.MM1_s
+ N_VDD_XI1.XI132.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI1.XI131.XI0.MM1 N_XI1.G8_XI1.XI131.XI0.MM1_d
+ N_XI1.XI131.NET6_XI1.XI131.XI0.MM1_g N_VDD_XI1.XI131.XI0.MM1_s
+ N_VDD_XI1.XI131.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI1.XI111.XI0.MM1 N_XI1.G7_XI1.XI111.XI0.MM1_d
+ N_XI1.XI111.NET6_XI1.XI111.XI0.MM1_g N_VDD_XI1.XI111.XI0.MM1_s
+ N_VDD_XI1.XI111.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI1.XI110.XI0.MM1 N_XI1.G6_XI1.XI110.XI0.MM1_d
+ N_XI1.XI110.NET6_XI1.XI110.XI0.MM1_g N_VDD_XI1.XI110.XI0.MM1_s
+ N_VDD_XI1.XI110.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI1.XI103.XI0.MM1 N_XI1.G5_XI1.XI103.XI0.MM1_d
+ N_XI1.XI103.NET6_XI1.XI103.XI0.MM1_g N_VDD_XI1.XI103.XI0.MM1_s
+ N_VDD_XI1.XI103.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI1.XI102.XI0.MM1 N_XI1.G4_XI1.XI102.XI0.MM1_d
+ N_XI1.XI102.NET6_XI1.XI102.XI0.MM1_g N_VDD_XI1.XI102.XI0.MM1_s
+ N_VDD_XI1.XI102.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI1.XI88.XI0.MM1 N_XI1.G3_XI1.XI88.XI0.MM1_d N_XI1.XI88.NET6_XI1.XI88.XI0.MM1_g
+ N_VDD_XI1.XI88.XI0.MM1_s N_VDD_XI1.XI88.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI1.XI82.XI0.MM1 N_XI1.G2_XI1.XI82.XI0.MM1_d N_XI1.XI82.NET6_XI1.XI82.XI0.MM1_g
+ N_VDD_XI1.XI82.XI0.MM1_s N_VDD_XI1.XI82.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI1.XI10.XI0.MM1 N_XI1.G1_XI1.XI10.XI0.MM1_d N_XI1.XI10.NET6_XI1.XI10.XI0.MM1_g
+ N_VDD_XI1.XI10.XI0.MM1_s N_VDD_XI1.XI10.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI1.XI134.MM4 N_XI1.P16_XI1.XI134.MM4_d N_MAX15_XI1.XI134.MM4_g
+ N_XI1.XI134.NET25_XI1.XI134.MM4_s N_VDD_XI1.XI134.XI9.MM1_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.425e-12 AS=6.7125e-13 PD=1.9e-06 PS=8.95e-07
mXI1.XI137.XI9.MM1 N_XI1.XI137.NET43_XI1.XI137.XI9.MM1_d
+ N_NET629_XI1.XI137.XI9.MM1_g N_VDD_XI1.XI137.XI9.MM1_s
+ N_VDD_XI1.XI153.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI1.XI140.XI9.MM1 N_XI1.XI140.NET43_XI1.XI140.XI9.MM1_d
+ N_NET630_XI1.XI140.XI9.MM1_g N_VDD_XI1.XI140.XI9.MM1_s
+ N_VDD_XI1.XI154.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI1.XI149.XI9.MM1 N_XI1.XI149.NET43_XI1.XI149.XI9.MM1_d
+ N_NET631_XI1.XI149.XI9.MM1_g N_VDD_XI1.XI149.XI9.MM1_s
+ N_VDD_XI1.XI157.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI1.XI146.XI9.MM1 N_XI1.XI146.NET43_XI1.XI146.XI9.MM1_d
+ N_NET632_XI1.XI146.XI9.MM1_g N_VDD_XI1.XI146.XI9.MM1_s
+ N_VDD_XI1.XI156.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI1.XI143.XI9.MM1 N_XI1.XI143.NET43_XI1.XI143.XI9.MM1_d
+ N_NET633_XI1.XI143.XI9.MM1_g N_VDD_XI1.XI143.XI9.MM1_s
+ N_VDD_XI1.XI155.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI1.XI128.XI9.MM1 N_XI1.XI128.NET43_XI1.XI128.XI9.MM1_d
+ N_NET634_XI1.XI128.XI9.MM1_g N_VDD_XI1.XI128.XI9.MM1_s
+ N_VDD_XI1.XI133.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI1.XI125.XI9.MM1 N_XI1.XI125.NET43_XI1.XI125.XI9.MM1_d
+ N_NET635_XI1.XI125.XI9.MM1_g N_VDD_XI1.XI125.XI9.MM1_s
+ N_VDD_XI1.XI132.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI1.XI122.XI9.MM1 N_XI1.XI122.NET43_XI1.XI122.XI9.MM1_d
+ N_NET636_XI1.XI122.XI9.MM1_g N_VDD_XI1.XI122.XI9.MM1_s
+ N_VDD_XI1.XI131.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI1.XI114.XI9.MM1 N_XI1.XI114.NET43_XI1.XI114.XI9.MM1_d
+ N_NET637_XI1.XI114.XI9.MM1_g N_VDD_XI1.XI114.XI9.MM1_s
+ N_VDD_XI1.XI111.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI1.XI109.XI9.MM1 N_XI1.XI109.NET43_XI1.XI109.XI9.MM1_d
+ N_NET638_XI1.XI109.XI9.MM1_g N_VDD_XI1.XI109.XI9.MM1_s
+ N_VDD_XI1.XI110.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI1.XI106.XI9.MM1 N_XI1.XI106.NET43_XI1.XI106.XI9.MM1_d
+ N_NET639_XI1.XI106.XI9.MM1_g N_VDD_XI1.XI106.XI9.MM1_s
+ N_VDD_XI1.XI103.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI1.XI101.XI9.MM1 N_XI1.XI101.NET43_XI1.XI101.XI9.MM1_d
+ N_NET640_XI1.XI101.XI9.MM1_g N_VDD_XI1.XI101.XI9.MM1_s
+ N_VDD_XI1.XI102.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI1.XI86.XI9.MM1 N_XI1.XI86.NET43_XI1.XI86.XI9.MM1_d
+ N_NET641_XI1.XI86.XI9.MM1_g N_VDD_XI1.XI86.XI9.MM1_s N_VDD_XI1.XI88.XI1.MM3_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI1.XI80.XI9.MM1 N_XI1.XI80.NET43_XI1.XI80.XI9.MM1_d
+ N_NET642_XI1.XI80.XI9.MM1_g N_VDD_XI1.XI80.XI9.MM1_s N_VDD_XI1.XI82.XI1.MM3_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI1.XI26.XI9.MM1 N_XI1.XI26.NET43_XI1.XI26.XI9.MM1_d
+ N_NET643_XI1.XI26.XI9.MM1_g N_VDD_XI1.XI26.XI9.MM1_s N_VDD_XI1.XI10.XI1.MM3_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI1.XI134.MM3 N_XI1.P16_XI1.XI134.MM3_d N_XI1.XI134.NET39_XI1.XI134.MM3_g
+ N_XI1.XI134.NET37_XI1.XI134.MM3_s N_VDD_XI1.XI134.XI9.MM1_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.425e-12 AS=5.4375e-13 PD=1.9e-06 PS=7.25e-07
mXI1.XI134.MM1 N_XI1.XI134.NET37_XI1.XI134.MM1_d N_NET628_XI1.XI134.MM1_g
+ N_VDD_XI1.XI134.MM1_s N_VDD_XI1.XI134.XI9.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=5.4375e-13 AS=7.65e-13 PD=7.25e-07 PS=2.52e-06
mXI1.XI137.MM5 N_XI1.XI137.NET25_XI1.XI137.MM5_d
+ N_XI1.XI137.NET43_XI1.XI137.MM5_g N_VDD_XI1.XI137.MM5_s
+ N_VDD_XI1.XI153.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=6.7125e-13 AS=9.675e-13
+ PD=8.95e-07 PS=2.79e-06
mXI1.XI140.MM5 N_XI1.XI140.NET25_XI1.XI140.MM5_d
+ N_XI1.XI140.NET43_XI1.XI140.MM5_g N_VDD_XI1.XI140.MM5_s
+ N_VDD_XI1.XI154.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=6.7125e-13 AS=9.675e-13
+ PD=8.95e-07 PS=2.79e-06
mXI1.XI149.MM5 N_XI1.XI149.NET25_XI1.XI149.MM5_d
+ N_XI1.XI149.NET43_XI1.XI149.MM5_g N_VDD_XI1.XI149.MM5_s
+ N_VDD_XI1.XI157.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=6.7125e-13 AS=9.675e-13
+ PD=8.95e-07 PS=2.79e-06
mXI1.XI146.MM5 N_XI1.XI146.NET25_XI1.XI146.MM5_d
+ N_XI1.XI146.NET43_XI1.XI146.MM5_g N_VDD_XI1.XI146.MM5_s
+ N_VDD_XI1.XI156.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=6.7125e-13 AS=9.675e-13
+ PD=8.95e-07 PS=2.79e-06
mXI1.XI143.MM5 N_XI1.XI143.NET25_XI1.XI143.MM5_d
+ N_XI1.XI143.NET43_XI1.XI143.MM5_g N_VDD_XI1.XI143.MM5_s
+ N_VDD_XI1.XI155.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=6.7125e-13 AS=9.675e-13
+ PD=8.95e-07 PS=2.79e-06
mXI1.XI128.MM5 N_XI1.XI128.NET25_XI1.XI128.MM5_d
+ N_XI1.XI128.NET43_XI1.XI128.MM5_g N_VDD_XI1.XI128.MM5_s
+ N_VDD_XI1.XI133.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=6.7125e-13 AS=9.675e-13
+ PD=8.95e-07 PS=2.79e-06
mXI1.XI125.MM5 N_XI1.XI125.NET25_XI1.XI125.MM5_d
+ N_XI1.XI125.NET43_XI1.XI125.MM5_g N_VDD_XI1.XI125.MM5_s
+ N_VDD_XI1.XI132.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=6.7125e-13 AS=9.675e-13
+ PD=8.95e-07 PS=2.79e-06
mXI1.XI122.MM5 N_XI1.XI122.NET25_XI1.XI122.MM5_d
+ N_XI1.XI122.NET43_XI1.XI122.MM5_g N_VDD_XI1.XI122.MM5_s
+ N_VDD_XI1.XI131.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=6.7125e-13 AS=9.675e-13
+ PD=8.95e-07 PS=2.79e-06
mXI1.XI114.MM5 N_XI1.XI114.NET25_XI1.XI114.MM5_d
+ N_XI1.XI114.NET43_XI1.XI114.MM5_g N_VDD_XI1.XI114.MM5_s
+ N_VDD_XI1.XI111.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=6.7125e-13 AS=9.675e-13
+ PD=8.95e-07 PS=2.79e-06
mXI1.XI109.MM5 N_XI1.XI109.NET25_XI1.XI109.MM5_d
+ N_XI1.XI109.NET43_XI1.XI109.MM5_g N_VDD_XI1.XI109.MM5_s
+ N_VDD_XI1.XI110.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=6.7125e-13 AS=9.675e-13
+ PD=8.95e-07 PS=2.79e-06
mXI1.XI106.MM5 N_XI1.XI106.NET25_XI1.XI106.MM5_d
+ N_XI1.XI106.NET43_XI1.XI106.MM5_g N_VDD_XI1.XI106.MM5_s
+ N_VDD_XI1.XI103.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=6.7125e-13 AS=9.675e-13
+ PD=8.95e-07 PS=2.79e-06
mXI1.XI101.MM5 N_XI1.XI101.NET25_XI1.XI101.MM5_d
+ N_XI1.XI101.NET43_XI1.XI101.MM5_g N_VDD_XI1.XI101.MM5_s
+ N_VDD_XI1.XI102.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=6.7125e-13 AS=9.675e-13
+ PD=8.95e-07 PS=2.79e-06
mXI1.XI86.MM5 N_XI1.XI86.NET25_XI1.XI86.MM5_d N_XI1.XI86.NET43_XI1.XI86.MM5_g
+ N_VDD_XI1.XI86.MM5_s N_VDD_XI1.XI88.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=6.7125e-13 AS=9.675e-13 PD=8.95e-07 PS=2.79e-06
mXI1.XI80.MM5 N_XI1.XI80.NET25_XI1.XI80.MM5_d N_XI1.XI80.NET43_XI1.XI80.MM5_g
+ N_VDD_XI1.XI80.MM5_s N_VDD_XI1.XI82.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=6.7125e-13 AS=9.675e-13 PD=8.95e-07 PS=2.79e-06
mXI1.XI26.MM5 N_XI1.XI26.NET25_XI1.XI26.MM5_d N_XI1.XI26.NET43_XI1.XI26.MM5_g
+ N_VDD_XI1.XI26.MM5_s N_VDD_XI1.XI10.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=6.7125e-13 AS=9.675e-13 PD=8.95e-07 PS=2.79e-06
mXI1.XI137.MM4 N_XI1.P15_XI1.XI137.MM4_d N_MAX14_XI1.XI137.MM4_g
+ N_XI1.XI137.NET25_XI1.XI137.MM4_s N_VDD_XI1.XI153.XI1.MM3_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.425e-12 AS=6.7125e-13 PD=1.9e-06 PS=8.95e-07
mXI1.XI140.MM4 N_XI1.P14_XI1.XI140.MM4_d N_MAX13_XI1.XI140.MM4_g
+ N_XI1.XI140.NET25_XI1.XI140.MM4_s N_VDD_XI1.XI154.XI1.MM3_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.425e-12 AS=6.7125e-13 PD=1.9e-06 PS=8.95e-07
mXI1.XI149.MM4 N_XI1.P13_XI1.XI149.MM4_d N_MAX12_XI1.XI149.MM4_g
+ N_XI1.XI149.NET25_XI1.XI149.MM4_s N_VDD_XI1.XI157.XI1.MM3_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.425e-12 AS=6.7125e-13 PD=1.9e-06 PS=8.95e-07
mXI1.XI146.MM4 N_XI1.P12_XI1.XI146.MM4_d N_MAX11_XI1.XI146.MM4_g
+ N_XI1.XI146.NET25_XI1.XI146.MM4_s N_VDD_XI1.XI156.XI1.MM3_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.425e-12 AS=6.7125e-13 PD=1.9e-06 PS=8.95e-07
mXI1.XI143.MM4 N_XI1.P11_XI1.XI143.MM4_d N_MAX10_XI1.XI143.MM4_g
+ N_XI1.XI143.NET25_XI1.XI143.MM4_s N_VDD_XI1.XI155.XI1.MM3_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.425e-12 AS=6.7125e-13 PD=1.9e-06 PS=8.95e-07
mXI1.XI128.MM4 N_XI1.P10_XI1.XI128.MM4_d N_MAX9_XI1.XI128.MM4_g
+ N_XI1.XI128.NET25_XI1.XI128.MM4_s N_VDD_XI1.XI133.XI1.MM3_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.425e-12 AS=6.7125e-13 PD=1.9e-06 PS=8.95e-07
mXI1.XI125.MM4 N_XI1.P9_XI1.XI125.MM4_d N_MAX8_XI1.XI125.MM4_g
+ N_XI1.XI125.NET25_XI1.XI125.MM4_s N_VDD_XI1.XI132.XI1.MM3_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.425e-12 AS=6.7125e-13 PD=1.9e-06 PS=8.95e-07
mXI1.XI122.MM4 N_XI1.P8_XI1.XI122.MM4_d N_MAX7_XI1.XI122.MM4_g
+ N_XI1.XI122.NET25_XI1.XI122.MM4_s N_VDD_XI1.XI131.XI1.MM3_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.425e-12 AS=6.7125e-13 PD=1.9e-06 PS=8.95e-07
mXI1.XI114.MM4 N_XI1.P7_XI1.XI114.MM4_d N_MAX6_XI1.XI114.MM4_g
+ N_XI1.XI114.NET25_XI1.XI114.MM4_s N_VDD_XI1.XI111.XI1.MM3_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.425e-12 AS=6.7125e-13 PD=1.9e-06 PS=8.95e-07
mXI1.XI109.MM4 N_XI1.P6_XI1.XI109.MM4_d N_MAX5_XI1.XI109.MM4_g
+ N_XI1.XI109.NET25_XI1.XI109.MM4_s N_VDD_XI1.XI110.XI1.MM3_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.425e-12 AS=6.7125e-13 PD=1.9e-06 PS=8.95e-07
mXI1.XI106.MM4 N_XI1.P5_XI1.XI106.MM4_d N_MAX4_XI1.XI106.MM4_g
+ N_XI1.XI106.NET25_XI1.XI106.MM4_s N_VDD_XI1.XI103.XI1.MM3_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.425e-12 AS=6.7125e-13 PD=1.9e-06 PS=8.95e-07
mXI1.XI101.MM4 N_XI1.P4_XI1.XI101.MM4_d N_MAX3_XI1.XI101.MM4_g
+ N_XI1.XI101.NET25_XI1.XI101.MM4_s N_VDD_XI1.XI102.XI1.MM3_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.425e-12 AS=6.7125e-13 PD=1.9e-06 PS=8.95e-07
mXI1.XI86.MM4 N_XI1.P3_XI1.XI86.MM4_d N_MAX2_XI1.XI86.MM4_g
+ N_XI1.XI86.NET25_XI1.XI86.MM4_s N_VDD_XI1.XI88.XI1.MM3_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.425e-12 AS=6.7125e-13 PD=1.9e-06 PS=8.95e-07
mXI1.XI80.MM4 N_XI1.P2_XI1.XI80.MM4_d N_MAX1_XI1.XI80.MM4_g
+ N_XI1.XI80.NET25_XI1.XI80.MM4_s N_VDD_XI1.XI82.XI1.MM3_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.425e-12 AS=6.7125e-13 PD=1.9e-06 PS=8.95e-07
mXI1.XI26.MM4 N_XI1.P1_XI1.XI26.MM4_d N_MAX0_XI1.XI26.MM4_g
+ N_XI1.XI26.NET25_XI1.XI26.MM4_s N_VDD_XI1.XI10.XI1.MM3_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.425e-12 AS=6.7125e-13 PD=1.9e-06 PS=8.95e-07
mXI1.XI134.XI4.MM1 N_XI1.XI134.NET39_XI1.XI134.XI4.MM1_d
+ N_MAX15_XI1.XI134.XI4.MM1_g N_VDD_XI1.XI134.XI4.MM1_s
+ N_VDD_XI1.XI134.XI9.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI1.XI137.MM3 N_XI1.P15_XI1.XI137.MM3_d N_XI1.XI137.NET39_XI1.XI137.MM3_g
+ N_XI1.XI137.NET37_XI1.XI137.MM3_s N_VDD_XI1.XI153.XI1.MM3_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.425e-12 AS=5.4375e-13 PD=1.9e-06 PS=7.25e-07
mXI1.XI140.MM3 N_XI1.P14_XI1.XI140.MM3_d N_XI1.XI140.NET39_XI1.XI140.MM3_g
+ N_XI1.XI140.NET37_XI1.XI140.MM3_s N_VDD_XI1.XI154.XI1.MM3_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.425e-12 AS=5.4375e-13 PD=1.9e-06 PS=7.25e-07
mXI1.XI149.MM3 N_XI1.P13_XI1.XI149.MM3_d N_XI1.XI149.NET39_XI1.XI149.MM3_g
+ N_XI1.XI149.NET37_XI1.XI149.MM3_s N_VDD_XI1.XI157.XI1.MM3_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.425e-12 AS=5.4375e-13 PD=1.9e-06 PS=7.25e-07
mXI1.XI146.MM3 N_XI1.P12_XI1.XI146.MM3_d N_XI1.XI146.NET39_XI1.XI146.MM3_g
+ N_XI1.XI146.NET37_XI1.XI146.MM3_s N_VDD_XI1.XI156.XI1.MM3_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.425e-12 AS=5.4375e-13 PD=1.9e-06 PS=7.25e-07
mXI1.XI143.MM3 N_XI1.P11_XI1.XI143.MM3_d N_XI1.XI143.NET39_XI1.XI143.MM3_g
+ N_XI1.XI143.NET37_XI1.XI143.MM3_s N_VDD_XI1.XI155.XI1.MM3_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.425e-12 AS=5.4375e-13 PD=1.9e-06 PS=7.25e-07
mXI1.XI128.MM3 N_XI1.P10_XI1.XI128.MM3_d N_XI1.XI128.NET39_XI1.XI128.MM3_g
+ N_XI1.XI128.NET37_XI1.XI128.MM3_s N_VDD_XI1.XI133.XI1.MM3_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.425e-12 AS=5.4375e-13 PD=1.9e-06 PS=7.25e-07
mXI1.XI125.MM3 N_XI1.P9_XI1.XI125.MM3_d N_XI1.XI125.NET39_XI1.XI125.MM3_g
+ N_XI1.XI125.NET37_XI1.XI125.MM3_s N_VDD_XI1.XI132.XI1.MM3_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.425e-12 AS=5.4375e-13 PD=1.9e-06 PS=7.25e-07
mXI1.XI122.MM3 N_XI1.P8_XI1.XI122.MM3_d N_XI1.XI122.NET39_XI1.XI122.MM3_g
+ N_XI1.XI122.NET37_XI1.XI122.MM3_s N_VDD_XI1.XI131.XI1.MM3_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.425e-12 AS=5.4375e-13 PD=1.9e-06 PS=7.25e-07
mXI1.XI114.MM3 N_XI1.P7_XI1.XI114.MM3_d N_XI1.XI114.NET39_XI1.XI114.MM3_g
+ N_XI1.XI114.NET37_XI1.XI114.MM3_s N_VDD_XI1.XI111.XI1.MM3_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.425e-12 AS=5.4375e-13 PD=1.9e-06 PS=7.25e-07
mXI1.XI109.MM3 N_XI1.P6_XI1.XI109.MM3_d N_XI1.XI109.NET39_XI1.XI109.MM3_g
+ N_XI1.XI109.NET37_XI1.XI109.MM3_s N_VDD_XI1.XI110.XI1.MM3_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.425e-12 AS=5.4375e-13 PD=1.9e-06 PS=7.25e-07
mXI1.XI106.MM3 N_XI1.P5_XI1.XI106.MM3_d N_XI1.XI106.NET39_XI1.XI106.MM3_g
+ N_XI1.XI106.NET37_XI1.XI106.MM3_s N_VDD_XI1.XI103.XI1.MM3_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.425e-12 AS=5.4375e-13 PD=1.9e-06 PS=7.25e-07
mXI1.XI101.MM3 N_XI1.P4_XI1.XI101.MM3_d N_XI1.XI101.NET39_XI1.XI101.MM3_g
+ N_XI1.XI101.NET37_XI1.XI101.MM3_s N_VDD_XI1.XI102.XI1.MM3_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.425e-12 AS=5.4375e-13 PD=1.9e-06 PS=7.25e-07
mXI1.XI86.MM3 N_XI1.P3_XI1.XI86.MM3_d N_XI1.XI86.NET39_XI1.XI86.MM3_g
+ N_XI1.XI86.NET37_XI1.XI86.MM3_s N_VDD_XI1.XI88.XI1.MM3_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.425e-12 AS=5.4375e-13 PD=1.9e-06 PS=7.25e-07
mXI1.XI80.MM3 N_XI1.P2_XI1.XI80.MM3_d N_XI1.XI80.NET39_XI1.XI80.MM3_g
+ N_XI1.XI80.NET37_XI1.XI80.MM3_s N_VDD_XI1.XI82.XI1.MM3_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.425e-12 AS=5.4375e-13 PD=1.9e-06 PS=7.25e-07
mXI1.XI26.MM3 N_XI1.P1_XI1.XI26.MM3_d N_XI1.XI26.NET39_XI1.XI26.MM3_g
+ N_XI1.XI26.NET37_XI1.XI26.MM3_s N_VDD_XI1.XI10.XI1.MM3_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.425e-12 AS=5.4375e-13 PD=1.9e-06 PS=7.25e-07
mXI1.XI137.MM1 N_XI1.XI137.NET37_XI1.XI137.MM1_d N_NET629_XI1.XI137.MM1_g
+ N_VDD_XI1.XI137.MM1_s N_VDD_XI1.XI153.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=5.4375e-13 AS=7.65e-13 PD=7.25e-07 PS=2.52e-06
mXI1.XI140.MM1 N_XI1.XI140.NET37_XI1.XI140.MM1_d N_NET630_XI1.XI140.MM1_g
+ N_VDD_XI1.XI140.MM1_s N_VDD_XI1.XI154.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=5.4375e-13 AS=7.65e-13 PD=7.25e-07 PS=2.52e-06
mXI1.XI149.MM1 N_XI1.XI149.NET37_XI1.XI149.MM1_d N_NET631_XI1.XI149.MM1_g
+ N_VDD_XI1.XI149.MM1_s N_VDD_XI1.XI157.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=5.4375e-13 AS=7.65e-13 PD=7.25e-07 PS=2.52e-06
mXI1.XI146.MM1 N_XI1.XI146.NET37_XI1.XI146.MM1_d N_NET632_XI1.XI146.MM1_g
+ N_VDD_XI1.XI146.MM1_s N_VDD_XI1.XI156.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=5.4375e-13 AS=7.65e-13 PD=7.25e-07 PS=2.52e-06
mXI1.XI143.MM1 N_XI1.XI143.NET37_XI1.XI143.MM1_d N_NET633_XI1.XI143.MM1_g
+ N_VDD_XI1.XI143.MM1_s N_VDD_XI1.XI155.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=5.4375e-13 AS=7.65e-13 PD=7.25e-07 PS=2.52e-06
mXI1.XI128.MM1 N_XI1.XI128.NET37_XI1.XI128.MM1_d N_NET634_XI1.XI128.MM1_g
+ N_VDD_XI1.XI128.MM1_s N_VDD_XI1.XI133.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=5.4375e-13 AS=7.65e-13 PD=7.25e-07 PS=2.52e-06
mXI1.XI125.MM1 N_XI1.XI125.NET37_XI1.XI125.MM1_d N_NET635_XI1.XI125.MM1_g
+ N_VDD_XI1.XI125.MM1_s N_VDD_XI1.XI132.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=5.4375e-13 AS=7.65e-13 PD=7.25e-07 PS=2.52e-06
mXI1.XI122.MM1 N_XI1.XI122.NET37_XI1.XI122.MM1_d N_NET636_XI1.XI122.MM1_g
+ N_VDD_XI1.XI122.MM1_s N_VDD_XI1.XI131.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=5.4375e-13 AS=7.65e-13 PD=7.25e-07 PS=2.52e-06
mXI1.XI114.MM1 N_XI1.XI114.NET37_XI1.XI114.MM1_d N_NET637_XI1.XI114.MM1_g
+ N_VDD_XI1.XI114.MM1_s N_VDD_XI1.XI111.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=5.4375e-13 AS=7.65e-13 PD=7.25e-07 PS=2.52e-06
mXI1.XI109.MM1 N_XI1.XI109.NET37_XI1.XI109.MM1_d N_NET638_XI1.XI109.MM1_g
+ N_VDD_XI1.XI109.MM1_s N_VDD_XI1.XI110.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=5.4375e-13 AS=7.65e-13 PD=7.25e-07 PS=2.52e-06
mXI1.XI106.MM1 N_XI1.XI106.NET37_XI1.XI106.MM1_d N_NET639_XI1.XI106.MM1_g
+ N_VDD_XI1.XI106.MM1_s N_VDD_XI1.XI103.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=5.4375e-13 AS=7.65e-13 PD=7.25e-07 PS=2.52e-06
mXI1.XI101.MM1 N_XI1.XI101.NET37_XI1.XI101.MM1_d N_NET640_XI1.XI101.MM1_g
+ N_VDD_XI1.XI101.MM1_s N_VDD_XI1.XI102.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=5.4375e-13 AS=7.65e-13 PD=7.25e-07 PS=2.52e-06
mXI1.XI86.MM1 N_XI1.XI86.NET37_XI1.XI86.MM1_d N_NET641_XI1.XI86.MM1_g
+ N_VDD_XI1.XI86.MM1_s N_VDD_XI1.XI88.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=5.4375e-13 AS=7.65e-13 PD=7.25e-07 PS=2.52e-06
mXI1.XI80.MM1 N_XI1.XI80.NET37_XI1.XI80.MM1_d N_NET642_XI1.XI80.MM1_g
+ N_VDD_XI1.XI80.MM1_s N_VDD_XI1.XI82.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=5.4375e-13 AS=7.65e-13 PD=7.25e-07 PS=2.52e-06
mXI1.XI26.MM1 N_XI1.XI26.NET37_XI1.XI26.MM1_d N_NET643_XI1.XI26.MM1_g
+ N_VDD_XI1.XI26.MM1_s N_VDD_XI1.XI10.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=5.4375e-13 AS=7.65e-13 PD=7.25e-07 PS=2.52e-06
mXI1.XI182.XI9.MM1 N_XI1.XI182.NET43_XI1.XI182.XI9.MM1_d
+ N_XI1.P16_XI1.XI182.XI9.MM1_g N_VDD_XI1.XI182.XI9.MM1_s
+ N_VDD_XI1.XI134.XI9.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI1.XI137.XI4.MM1 N_XI1.XI137.NET39_XI1.XI137.XI4.MM1_d
+ N_MAX14_XI1.XI137.XI4.MM1_g N_VDD_XI1.XI137.XI4.MM1_s
+ N_VDD_XI1.XI153.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI1.XI140.XI4.MM1 N_XI1.XI140.NET39_XI1.XI140.XI4.MM1_d
+ N_MAX13_XI1.XI140.XI4.MM1_g N_VDD_XI1.XI140.XI4.MM1_s
+ N_VDD_XI1.XI154.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI1.XI149.XI4.MM1 N_XI1.XI149.NET39_XI1.XI149.XI4.MM1_d
+ N_MAX12_XI1.XI149.XI4.MM1_g N_VDD_XI1.XI149.XI4.MM1_s
+ N_VDD_XI1.XI157.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI1.XI146.XI4.MM1 N_XI1.XI146.NET39_XI1.XI146.XI4.MM1_d
+ N_MAX11_XI1.XI146.XI4.MM1_g N_VDD_XI1.XI146.XI4.MM1_s
+ N_VDD_XI1.XI156.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI1.XI143.XI4.MM1 N_XI1.XI143.NET39_XI1.XI143.XI4.MM1_d
+ N_MAX10_XI1.XI143.XI4.MM1_g N_VDD_XI1.XI143.XI4.MM1_s
+ N_VDD_XI1.XI155.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI1.XI128.XI4.MM1 N_XI1.XI128.NET39_XI1.XI128.XI4.MM1_d
+ N_MAX9_XI1.XI128.XI4.MM1_g N_VDD_XI1.XI128.XI4.MM1_s N_VDD_XI1.XI133.XI1.MM3_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI1.XI125.XI4.MM1 N_XI1.XI125.NET39_XI1.XI125.XI4.MM1_d
+ N_MAX8_XI1.XI125.XI4.MM1_g N_VDD_XI1.XI125.XI4.MM1_s N_VDD_XI1.XI132.XI1.MM3_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI1.XI122.XI4.MM1 N_XI1.XI122.NET39_XI1.XI122.XI4.MM1_d
+ N_MAX7_XI1.XI122.XI4.MM1_g N_VDD_XI1.XI122.XI4.MM1_s N_VDD_XI1.XI131.XI1.MM3_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI1.XI114.XI4.MM1 N_XI1.XI114.NET39_XI1.XI114.XI4.MM1_d
+ N_MAX6_XI1.XI114.XI4.MM1_g N_VDD_XI1.XI114.XI4.MM1_s N_VDD_XI1.XI111.XI1.MM3_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI1.XI109.XI4.MM1 N_XI1.XI109.NET39_XI1.XI109.XI4.MM1_d
+ N_MAX5_XI1.XI109.XI4.MM1_g N_VDD_XI1.XI109.XI4.MM1_s N_VDD_XI1.XI110.XI1.MM3_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI1.XI106.XI4.MM1 N_XI1.XI106.NET39_XI1.XI106.XI4.MM1_d
+ N_MAX4_XI1.XI106.XI4.MM1_g N_VDD_XI1.XI106.XI4.MM1_s N_VDD_XI1.XI103.XI1.MM3_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI1.XI101.XI4.MM1 N_XI1.XI101.NET39_XI1.XI101.XI4.MM1_d
+ N_MAX3_XI1.XI101.XI4.MM1_g N_VDD_XI1.XI101.XI4.MM1_s N_VDD_XI1.XI102.XI1.MM3_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI1.XI86.XI4.MM1 N_XI1.XI86.NET39_XI1.XI86.XI4.MM1_d N_MAX2_XI1.XI86.XI4.MM1_g
+ N_VDD_XI1.XI86.XI4.MM1_s N_VDD_XI1.XI88.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI1.XI80.XI4.MM1 N_XI1.XI80.NET39_XI1.XI80.XI4.MM1_d N_MAX1_XI1.XI80.XI4.MM1_g
+ N_VDD_XI1.XI80.XI4.MM1_s N_VDD_XI1.XI82.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI1.XI26.XI4.MM1 N_XI1.XI26.NET39_XI1.XI26.XI4.MM1_d N_MAX0_XI1.XI26.XI4.MM1_g
+ N_VDD_XI1.XI26.XI4.MM1_s N_VDD_XI1.XI10.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI1.XI182.MM5 N_XI1.XI182.NET25_XI1.XI182.MM5_d
+ N_XI1.XI182.NET43_XI1.XI182.MM5_g N_VDD_XI1.XI182.MM5_s
+ N_VDD_XI1.XI134.XI9.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=6.7125e-13 AS=9.675e-13
+ PD=8.95e-07 PS=2.79e-06
mXI1.XI168.XI1.XI1.MM1 N_XI1.XI168.XI1.NET6_XI1.XI168.XI1.XI1.MM1_d
+ N_XI1.NET288_XI1.XI168.XI1.XI1.MM1_g N_VDD_XI1.XI168.XI1.XI1.MM1_s
+ N_VDD_XI1.XI153.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.35e-13
+ PD=7.4e-07 PS=2.48e-06
mXI1.XI167.XI1.XI1.MM1 N_XI1.XI167.XI1.NET6_XI1.XI167.XI1.XI1.MM1_d
+ N_XI1.NET282_XI1.XI167.XI1.XI1.MM1_g N_VDD_XI1.XI167.XI1.XI1.MM1_s
+ N_VDD_XI1.XI154.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.35e-13
+ PD=7.4e-07 PS=2.48e-06
mXI1.XI166.XI1.XI1.MM1 N_XI1.XI166.XI1.NET6_XI1.XI166.XI1.XI1.MM1_d
+ N_XI1.NET276_XI1.XI166.XI1.XI1.MM1_g N_VDD_XI1.XI166.XI1.XI1.MM1_s
+ N_VDD_XI1.XI157.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.35e-13
+ PD=7.4e-07 PS=2.48e-06
mXI1.XI165.XI1.XI1.MM1 N_XI1.XI165.XI1.NET6_XI1.XI165.XI1.XI1.MM1_d
+ N_XI1.NET270_XI1.XI165.XI1.XI1.MM1_g N_VDD_XI1.XI165.XI1.XI1.MM1_s
+ N_VDD_XI1.XI156.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.35e-13
+ PD=7.4e-07 PS=2.48e-06
mXI1.XI159.XI1.XI1.MM1 N_XI1.XI159.XI1.NET6_XI1.XI159.XI1.XI1.MM1_d
+ N_XI1.NET246_XI1.XI159.XI1.XI1.MM1_g N_VDD_XI1.XI159.XI1.XI1.MM1_s
+ N_VDD_XI1.XI155.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.35e-13
+ PD=7.4e-07 PS=2.48e-06
mXI1.XI160.XI1.XI1.MM1 N_XI1.XI160.XI1.NET6_XI1.XI160.XI1.XI1.MM1_d
+ N_XI1.NET252_XI1.XI160.XI1.XI1.MM1_g N_VDD_XI1.XI160.XI1.XI1.MM1_s
+ N_VDD_XI1.XI133.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.35e-13
+ PD=7.4e-07 PS=2.48e-06
mXI1.XI161.XI1.XI1.MM1 N_XI1.XI161.XI1.NET6_XI1.XI161.XI1.XI1.MM1_d
+ N_XI1.NET258_XI1.XI161.XI1.XI1.MM1_g N_VDD_XI1.XI161.XI1.XI1.MM1_s
+ N_VDD_XI1.XI132.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.35e-13
+ PD=7.4e-07 PS=2.48e-06
mXI1.XI162.XI1.XI1.MM1 N_XI1.XI162.XI1.NET6_XI1.XI162.XI1.XI1.MM1_d
+ N_XI1.NET264_XI1.XI162.XI1.XI1.MM1_g N_VDD_XI1.XI162.XI1.XI1.MM1_s
+ N_VDD_XI1.XI131.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.35e-13
+ PD=7.4e-07 PS=2.48e-06
mXI1.XI121.XI1.XI1.MM1 N_XI1.XI121.XI1.NET6_XI1.XI121.XI1.XI1.MM1_d
+ N_XI1.NET204_XI1.XI121.XI1.XI1.MM1_g N_VDD_XI1.XI121.XI1.XI1.MM1_s
+ N_VDD_XI1.XI111.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.35e-13
+ PD=7.4e-07 PS=2.48e-06
mXI1.XI120.XI1.XI1.MM1 N_XI1.XI120.XI1.NET6_XI1.XI120.XI1.XI1.MM1_d
+ N_XI1.NET210_XI1.XI120.XI1.XI1.MM1_g N_VDD_XI1.XI120.XI1.XI1.MM1_s
+ N_VDD_XI1.XI110.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.35e-13
+ PD=7.4e-07 PS=2.48e-06
mXI1.XI119.XI1.XI1.MM1 N_XI1.XI119.XI1.NET6_XI1.XI119.XI1.XI1.MM1_d
+ N_XI1.NET216_XI1.XI119.XI1.XI1.MM1_g N_VDD_XI1.XI119.XI1.XI1.MM1_s
+ N_VDD_XI1.XI103.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.35e-13
+ PD=7.4e-07 PS=2.48e-06
mXI1.XI118.XI1.XI1.MM1 N_XI1.XI118.XI1.NET6_XI1.XI118.XI1.XI1.MM1_d
+ N_XI1.NET222_XI1.XI118.XI1.XI1.MM1_g N_VDD_XI1.XI118.XI1.XI1.MM1_s
+ N_VDD_XI1.XI102.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.35e-13
+ PD=7.4e-07 PS=2.48e-06
mXI1.XI91.XI1.XI1.MM1 N_XI1.XI91.XI1.NET6_XI1.XI91.XI1.XI1.MM1_d
+ N_XI1.NET228_XI1.XI91.XI1.XI1.MM1_g N_VDD_XI1.XI91.XI1.XI1.MM1_s
+ N_VDD_XI1.XI88.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.35e-13
+ PD=7.4e-07 PS=2.48e-06
mXI1.XI90.XI1.XI1.MM1 N_XI1.XI90.XI1.NET6_XI1.XI90.XI1.XI1.MM1_d
+ N_XI1.NET240_XI1.XI90.XI1.XI1.MM1_g N_VDD_XI1.XI90.XI1.XI1.MM1_s
+ N_VDD_XI1.XI82.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.35e-13
+ PD=7.4e-07 PS=2.48e-06
mXI1.XI89.XI1.XI1.MM1 N_XI1.XI89.XI1.NET6_XI1.XI89.XI1.XI1.MM1_d
+ N_CIN2_XI1.XI89.XI1.XI1.MM1_g N_VDD_XI1.XI89.XI1.XI1.MM1_s
+ N_VDD_XI1.XI10.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.35e-13
+ PD=7.4e-07 PS=2.48e-06
mXI1.XI182.MM4 N_NET105_XI1.XI182.MM4_d N_XI1.NET198_XI1.XI182.MM4_g
+ N_XI1.XI182.NET25_XI1.XI182.MM4_s N_VDD_XI1.XI134.XI9.MM1_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.425e-12 AS=6.7125e-13 PD=1.9e-06 PS=8.95e-07
mXI1.XI168.XI1.XI1.MM3 N_XI1.XI168.XI1.NET6_XI1.XI168.XI1.XI1.MM3_d
+ N_XI1.P15_XI1.XI168.XI1.XI1.MM3_g N_VDD_XI1.XI168.XI1.XI1.MM3_s
+ N_VDD_XI1.XI153.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.65e-13
+ PD=7.4e-07 PS=2.52e-06
mXI1.XI167.XI1.XI1.MM3 N_XI1.XI167.XI1.NET6_XI1.XI167.XI1.XI1.MM3_d
+ N_XI1.P14_XI1.XI167.XI1.XI1.MM3_g N_VDD_XI1.XI167.XI1.XI1.MM3_s
+ N_VDD_XI1.XI154.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.65e-13
+ PD=7.4e-07 PS=2.52e-06
mXI1.XI166.XI1.XI1.MM3 N_XI1.XI166.XI1.NET6_XI1.XI166.XI1.XI1.MM3_d
+ N_XI1.P13_XI1.XI166.XI1.XI1.MM3_g N_VDD_XI1.XI166.XI1.XI1.MM3_s
+ N_VDD_XI1.XI157.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.65e-13
+ PD=7.4e-07 PS=2.52e-06
mXI1.XI165.XI1.XI1.MM3 N_XI1.XI165.XI1.NET6_XI1.XI165.XI1.XI1.MM3_d
+ N_XI1.P12_XI1.XI165.XI1.XI1.MM3_g N_VDD_XI1.XI165.XI1.XI1.MM3_s
+ N_VDD_XI1.XI156.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.65e-13
+ PD=7.4e-07 PS=2.52e-06
mXI1.XI159.XI1.XI1.MM3 N_XI1.XI159.XI1.NET6_XI1.XI159.XI1.XI1.MM3_d
+ N_XI1.P11_XI1.XI159.XI1.XI1.MM3_g N_VDD_XI1.XI159.XI1.XI1.MM3_s
+ N_VDD_XI1.XI155.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.65e-13
+ PD=7.4e-07 PS=2.52e-06
mXI1.XI160.XI1.XI1.MM3 N_XI1.XI160.XI1.NET6_XI1.XI160.XI1.XI1.MM3_d
+ N_XI1.P10_XI1.XI160.XI1.XI1.MM3_g N_VDD_XI1.XI160.XI1.XI1.MM3_s
+ N_VDD_XI1.XI133.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.65e-13
+ PD=7.4e-07 PS=2.52e-06
mXI1.XI161.XI1.XI1.MM3 N_XI1.XI161.XI1.NET6_XI1.XI161.XI1.XI1.MM3_d
+ N_XI1.P9_XI1.XI161.XI1.XI1.MM3_g N_VDD_XI1.XI161.XI1.XI1.MM3_s
+ N_VDD_XI1.XI132.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.65e-13
+ PD=7.4e-07 PS=2.52e-06
mXI1.XI162.XI1.XI1.MM3 N_XI1.XI162.XI1.NET6_XI1.XI162.XI1.XI1.MM3_d
+ N_XI1.P8_XI1.XI162.XI1.XI1.MM3_g N_VDD_XI1.XI162.XI1.XI1.MM3_s
+ N_VDD_XI1.XI131.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.65e-13
+ PD=7.4e-07 PS=2.52e-06
mXI1.XI121.XI1.XI1.MM3 N_XI1.XI121.XI1.NET6_XI1.XI121.XI1.XI1.MM3_d
+ N_XI1.P7_XI1.XI121.XI1.XI1.MM3_g N_VDD_XI1.XI121.XI1.XI1.MM3_s
+ N_VDD_XI1.XI111.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.65e-13
+ PD=7.4e-07 PS=2.52e-06
mXI1.XI120.XI1.XI1.MM3 N_XI1.XI120.XI1.NET6_XI1.XI120.XI1.XI1.MM3_d
+ N_XI1.P6_XI1.XI120.XI1.XI1.MM3_g N_VDD_XI1.XI120.XI1.XI1.MM3_s
+ N_VDD_XI1.XI110.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.65e-13
+ PD=7.4e-07 PS=2.52e-06
mXI1.XI119.XI1.XI1.MM3 N_XI1.XI119.XI1.NET6_XI1.XI119.XI1.XI1.MM3_d
+ N_XI1.P5_XI1.XI119.XI1.XI1.MM3_g N_VDD_XI1.XI119.XI1.XI1.MM3_s
+ N_VDD_XI1.XI103.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.65e-13
+ PD=7.4e-07 PS=2.52e-06
mXI1.XI118.XI1.XI1.MM3 N_XI1.XI118.XI1.NET6_XI1.XI118.XI1.XI1.MM3_d
+ N_XI1.P4_XI1.XI118.XI1.XI1.MM3_g N_VDD_XI1.XI118.XI1.XI1.MM3_s
+ N_VDD_XI1.XI102.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.65e-13
+ PD=7.4e-07 PS=2.52e-06
mXI1.XI91.XI1.XI1.MM3 N_XI1.XI91.XI1.NET6_XI1.XI91.XI1.XI1.MM3_d
+ N_XI1.P3_XI1.XI91.XI1.XI1.MM3_g N_VDD_XI1.XI91.XI1.XI1.MM3_s
+ N_VDD_XI1.XI88.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.65e-13
+ PD=7.4e-07 PS=2.52e-06
mXI1.XI90.XI1.XI1.MM3 N_XI1.XI90.XI1.NET6_XI1.XI90.XI1.XI1.MM3_d
+ N_XI1.P2_XI1.XI90.XI1.XI1.MM3_g N_VDD_XI1.XI90.XI1.XI1.MM3_s
+ N_VDD_XI1.XI82.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.65e-13
+ PD=7.4e-07 PS=2.52e-06
mXI1.XI89.XI1.XI1.MM3 N_XI1.XI89.XI1.NET6_XI1.XI89.XI1.XI1.MM3_d
+ N_XI1.P1_XI1.XI89.XI1.XI1.MM3_g N_VDD_XI1.XI89.XI1.XI1.MM3_s
+ N_VDD_XI1.XI10.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=5.55e-13 AS=7.65e-13
+ PD=7.4e-07 PS=2.52e-06
mXI7.MM1 N_NET0855_XI7.MM1_d N_NET105_XI7.MM1_g N_VDD_XI7.MM1_s N_VDD_XI7.MM1_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI1.XI182.MM3 N_NET105_XI1.XI182.MM3_d N_XI1.XI182.NET39_XI1.XI182.MM3_g
+ N_XI1.XI182.NET37_XI1.XI182.MM3_s N_VDD_XI1.XI134.XI9.MM1_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.425e-12 AS=5.4375e-13 PD=1.9e-06 PS=7.25e-07
mXI1.XI168.XI1.XI0.MM1 N_XI1.XI168.NET13_XI1.XI168.XI1.XI0.MM1_d
+ N_XI1.XI168.XI1.NET6_XI1.XI168.XI1.XI0.MM1_g N_VDD_XI1.XI168.XI1.XI0.MM1_s
+ N_VDD_XI1.XI153.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI1.XI167.XI1.XI0.MM1 N_XI1.XI167.NET13_XI1.XI167.XI1.XI0.MM1_d
+ N_XI1.XI167.XI1.NET6_XI1.XI167.XI1.XI0.MM1_g N_VDD_XI1.XI167.XI1.XI0.MM1_s
+ N_VDD_XI1.XI154.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI1.XI166.XI1.XI0.MM1 N_XI1.XI166.NET13_XI1.XI166.XI1.XI0.MM1_d
+ N_XI1.XI166.XI1.NET6_XI1.XI166.XI1.XI0.MM1_g N_VDD_XI1.XI166.XI1.XI0.MM1_s
+ N_VDD_XI1.XI157.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI1.XI165.XI1.XI0.MM1 N_XI1.XI165.NET13_XI1.XI165.XI1.XI0.MM1_d
+ N_XI1.XI165.XI1.NET6_XI1.XI165.XI1.XI0.MM1_g N_VDD_XI1.XI165.XI1.XI0.MM1_s
+ N_VDD_XI1.XI156.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI1.XI159.XI1.XI0.MM1 N_XI1.XI159.NET13_XI1.XI159.XI1.XI0.MM1_d
+ N_XI1.XI159.XI1.NET6_XI1.XI159.XI1.XI0.MM1_g N_VDD_XI1.XI159.XI1.XI0.MM1_s
+ N_VDD_XI1.XI155.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI1.XI160.XI1.XI0.MM1 N_XI1.XI160.NET13_XI1.XI160.XI1.XI0.MM1_d
+ N_XI1.XI160.XI1.NET6_XI1.XI160.XI1.XI0.MM1_g N_VDD_XI1.XI160.XI1.XI0.MM1_s
+ N_VDD_XI1.XI133.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI1.XI161.XI1.XI0.MM1 N_XI1.XI161.NET13_XI1.XI161.XI1.XI0.MM1_d
+ N_XI1.XI161.XI1.NET6_XI1.XI161.XI1.XI0.MM1_g N_VDD_XI1.XI161.XI1.XI0.MM1_s
+ N_VDD_XI1.XI132.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI1.XI162.XI1.XI0.MM1 N_XI1.XI162.NET13_XI1.XI162.XI1.XI0.MM1_d
+ N_XI1.XI162.XI1.NET6_XI1.XI162.XI1.XI0.MM1_g N_VDD_XI1.XI162.XI1.XI0.MM1_s
+ N_VDD_XI1.XI131.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI1.XI121.XI1.XI0.MM1 N_XI1.XI121.NET13_XI1.XI121.XI1.XI0.MM1_d
+ N_XI1.XI121.XI1.NET6_XI1.XI121.XI1.XI0.MM1_g N_VDD_XI1.XI121.XI1.XI0.MM1_s
+ N_VDD_XI1.XI111.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI1.XI120.XI1.XI0.MM1 N_XI1.XI120.NET13_XI1.XI120.XI1.XI0.MM1_d
+ N_XI1.XI120.XI1.NET6_XI1.XI120.XI1.XI0.MM1_g N_VDD_XI1.XI120.XI1.XI0.MM1_s
+ N_VDD_XI1.XI110.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI1.XI119.XI1.XI0.MM1 N_XI1.XI119.NET13_XI1.XI119.XI1.XI0.MM1_d
+ N_XI1.XI119.XI1.NET6_XI1.XI119.XI1.XI0.MM1_g N_VDD_XI1.XI119.XI1.XI0.MM1_s
+ N_VDD_XI1.XI103.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI1.XI118.XI1.XI0.MM1 N_XI1.XI118.NET13_XI1.XI118.XI1.XI0.MM1_d
+ N_XI1.XI118.XI1.NET6_XI1.XI118.XI1.XI0.MM1_g N_VDD_XI1.XI118.XI1.XI0.MM1_s
+ N_VDD_XI1.XI102.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI1.XI91.XI1.XI0.MM1 N_XI1.XI91.NET13_XI1.XI91.XI1.XI0.MM1_d
+ N_XI1.XI91.XI1.NET6_XI1.XI91.XI1.XI0.MM1_g N_VDD_XI1.XI91.XI1.XI0.MM1_s
+ N_VDD_XI1.XI88.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI1.XI90.XI1.XI0.MM1 N_XI1.XI90.NET13_XI1.XI90.XI1.XI0.MM1_d
+ N_XI1.XI90.XI1.NET6_XI1.XI90.XI1.XI0.MM1_g N_VDD_XI1.XI90.XI1.XI0.MM1_s
+ N_VDD_XI1.XI82.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI1.XI89.XI1.XI0.MM1 N_XI1.XI89.NET13_XI1.XI89.XI1.XI0.MM1_d
+ N_XI1.XI89.XI1.NET6_XI1.XI89.XI1.XI0.MM1_g N_VDD_XI1.XI89.XI1.XI0.MM1_s
+ N_VDD_XI1.XI10.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI1.XI182.MM1 N_XI1.XI182.NET37_XI1.XI182.MM1_d N_XI1.P16_XI1.XI182.MM1_g
+ N_VDD_XI1.XI182.MM1_s N_VDD_XI1.XI134.XI9.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=5.4375e-13 AS=7.65e-13 PD=7.25e-07 PS=2.52e-06
mXI1.XI168.XI0.XI0.MM1 N_XI1.XI168.XI0.XI0.NET17_XI1.XI168.XI0.XI0.MM1_d
+ N_XI1.XI168.NET13_XI1.XI168.XI0.XI0.MM1_g N_VDD_XI1.XI168.XI0.XI0.MM1_s
+ N_VDD_XI1.XI153.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=4.125e-13 AS=7.35e-13
+ PD=5.5e-07 PS=2.48e-06
mXI1.XI167.XI0.XI0.MM1 N_XI1.XI167.XI0.XI0.NET17_XI1.XI167.XI0.XI0.MM1_d
+ N_XI1.XI167.NET13_XI1.XI167.XI0.XI0.MM1_g N_VDD_XI1.XI167.XI0.XI0.MM1_s
+ N_VDD_XI1.XI154.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=4.125e-13 AS=7.35e-13
+ PD=5.5e-07 PS=2.48e-06
mXI1.XI166.XI0.XI0.MM1 N_XI1.XI166.XI0.XI0.NET17_XI1.XI166.XI0.XI0.MM1_d
+ N_XI1.XI166.NET13_XI1.XI166.XI0.XI0.MM1_g N_VDD_XI1.XI166.XI0.XI0.MM1_s
+ N_VDD_XI1.XI157.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=4.125e-13 AS=7.35e-13
+ PD=5.5e-07 PS=2.48e-06
mXI1.XI165.XI0.XI0.MM1 N_XI1.XI165.XI0.XI0.NET17_XI1.XI165.XI0.XI0.MM1_d
+ N_XI1.XI165.NET13_XI1.XI165.XI0.XI0.MM1_g N_VDD_XI1.XI165.XI0.XI0.MM1_s
+ N_VDD_XI1.XI156.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=4.125e-13 AS=7.35e-13
+ PD=5.5e-07 PS=2.48e-06
mXI1.XI159.XI0.XI0.MM1 N_XI1.XI159.XI0.XI0.NET17_XI1.XI159.XI0.XI0.MM1_d
+ N_XI1.XI159.NET13_XI1.XI159.XI0.XI0.MM1_g N_VDD_XI1.XI159.XI0.XI0.MM1_s
+ N_VDD_XI1.XI155.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=4.125e-13 AS=7.35e-13
+ PD=5.5e-07 PS=2.48e-06
mXI1.XI160.XI0.XI0.MM1 N_XI1.XI160.XI0.XI0.NET17_XI1.XI160.XI0.XI0.MM1_d
+ N_XI1.XI160.NET13_XI1.XI160.XI0.XI0.MM1_g N_VDD_XI1.XI160.XI0.XI0.MM1_s
+ N_VDD_XI1.XI133.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=4.125e-13 AS=7.35e-13
+ PD=5.5e-07 PS=2.48e-06
mXI1.XI161.XI0.XI0.MM1 N_XI1.XI161.XI0.XI0.NET17_XI1.XI161.XI0.XI0.MM1_d
+ N_XI1.XI161.NET13_XI1.XI161.XI0.XI0.MM1_g N_VDD_XI1.XI161.XI0.XI0.MM1_s
+ N_VDD_XI1.XI132.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=4.125e-13 AS=7.35e-13
+ PD=5.5e-07 PS=2.48e-06
mXI1.XI162.XI0.XI0.MM1 N_XI1.XI162.XI0.XI0.NET17_XI1.XI162.XI0.XI0.MM1_d
+ N_XI1.XI162.NET13_XI1.XI162.XI0.XI0.MM1_g N_VDD_XI1.XI162.XI0.XI0.MM1_s
+ N_VDD_XI1.XI131.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=4.125e-13 AS=7.35e-13
+ PD=5.5e-07 PS=2.48e-06
mXI1.XI121.XI0.XI0.MM1 N_XI1.XI121.XI0.XI0.NET17_XI1.XI121.XI0.XI0.MM1_d
+ N_XI1.XI121.NET13_XI1.XI121.XI0.XI0.MM1_g N_VDD_XI1.XI121.XI0.XI0.MM1_s
+ N_VDD_XI1.XI111.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=4.125e-13 AS=7.35e-13
+ PD=5.5e-07 PS=2.48e-06
mXI1.XI120.XI0.XI0.MM1 N_XI1.XI120.XI0.XI0.NET17_XI1.XI120.XI0.XI0.MM1_d
+ N_XI1.XI120.NET13_XI1.XI120.XI0.XI0.MM1_g N_VDD_XI1.XI120.XI0.XI0.MM1_s
+ N_VDD_XI1.XI110.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=4.125e-13 AS=7.35e-13
+ PD=5.5e-07 PS=2.48e-06
mXI1.XI119.XI0.XI0.MM1 N_XI1.XI119.XI0.XI0.NET17_XI1.XI119.XI0.XI0.MM1_d
+ N_XI1.XI119.NET13_XI1.XI119.XI0.XI0.MM1_g N_VDD_XI1.XI119.XI0.XI0.MM1_s
+ N_VDD_XI1.XI103.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=4.125e-13 AS=7.35e-13
+ PD=5.5e-07 PS=2.48e-06
mXI1.XI118.XI0.XI0.MM1 N_XI1.XI118.XI0.XI0.NET17_XI1.XI118.XI0.XI0.MM1_d
+ N_XI1.XI118.NET13_XI1.XI118.XI0.XI0.MM1_g N_VDD_XI1.XI118.XI0.XI0.MM1_s
+ N_VDD_XI1.XI102.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=4.125e-13 AS=7.35e-13
+ PD=5.5e-07 PS=2.48e-06
mXI1.XI91.XI0.XI0.MM1 N_XI1.XI91.XI0.XI0.NET17_XI1.XI91.XI0.XI0.MM1_d
+ N_XI1.XI91.NET13_XI1.XI91.XI0.XI0.MM1_g N_VDD_XI1.XI91.XI0.XI0.MM1_s
+ N_VDD_XI1.XI88.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=4.125e-13 AS=7.35e-13
+ PD=5.5e-07 PS=2.48e-06
mXI1.XI90.XI0.XI0.MM1 N_XI1.XI90.XI0.XI0.NET17_XI1.XI90.XI0.XI0.MM1_d
+ N_XI1.XI90.NET13_XI1.XI90.XI0.XI0.MM1_g N_VDD_XI1.XI90.XI0.XI0.MM1_s
+ N_VDD_XI1.XI82.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=4.125e-13 AS=7.35e-13
+ PD=5.5e-07 PS=2.48e-06
mXI1.XI89.XI0.XI0.MM1 N_XI1.XI89.XI0.XI0.NET17_XI1.XI89.XI0.XI0.MM1_d
+ N_XI1.XI89.NET13_XI1.XI89.XI0.XI0.MM1_g N_VDD_XI1.XI89.XI0.XI0.MM1_s
+ N_VDD_XI1.XI10.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=4.125e-13 AS=7.35e-13
+ PD=5.5e-07 PS=2.48e-06
mXI1.XI182.XI4.MM1 N_XI1.XI182.NET39_XI1.XI182.XI4.MM1_d
+ N_XI1.NET198_XI1.XI182.XI4.MM1_g N_VDD_XI1.XI182.XI4.MM1_s
+ N_VDD_XI1.XI134.XI9.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI1.XI168.XI0.XI0.MM3 N_XI1.XI168.XI0.NET12_XI1.XI168.XI0.XI0.MM3_d
+ N_XI1.G15_XI1.XI168.XI0.XI0.MM3_g
+ N_XI1.XI168.XI0.XI0.NET17_XI1.XI168.XI0.XI0.MM3_s N_VDD_XI1.XI153.XI1.MM3_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=4.125e-13 PD=2.52e-06 PS=5.5e-07
mXI1.XI167.XI0.XI0.MM3 N_XI1.XI167.XI0.NET12_XI1.XI167.XI0.XI0.MM3_d
+ N_XI1.G14_XI1.XI167.XI0.XI0.MM3_g
+ N_XI1.XI167.XI0.XI0.NET17_XI1.XI167.XI0.XI0.MM3_s N_VDD_XI1.XI154.XI1.MM3_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=4.125e-13 PD=2.52e-06 PS=5.5e-07
mXI1.XI166.XI0.XI0.MM3 N_XI1.XI166.XI0.NET12_XI1.XI166.XI0.XI0.MM3_d
+ N_XI1.G13_XI1.XI166.XI0.XI0.MM3_g
+ N_XI1.XI166.XI0.XI0.NET17_XI1.XI166.XI0.XI0.MM3_s N_VDD_XI1.XI157.XI1.MM3_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=4.125e-13 PD=2.52e-06 PS=5.5e-07
mXI1.XI165.XI0.XI0.MM3 N_XI1.XI165.XI0.NET12_XI1.XI165.XI0.XI0.MM3_d
+ N_XI1.G12_XI1.XI165.XI0.XI0.MM3_g
+ N_XI1.XI165.XI0.XI0.NET17_XI1.XI165.XI0.XI0.MM3_s N_VDD_XI1.XI156.XI1.MM3_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=4.125e-13 PD=2.52e-06 PS=5.5e-07
mXI1.XI159.XI0.XI0.MM3 N_XI1.XI159.XI0.NET12_XI1.XI159.XI0.XI0.MM3_d
+ N_XI1.G11_XI1.XI159.XI0.XI0.MM3_g
+ N_XI1.XI159.XI0.XI0.NET17_XI1.XI159.XI0.XI0.MM3_s N_VDD_XI1.XI155.XI1.MM3_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=4.125e-13 PD=2.52e-06 PS=5.5e-07
mXI1.XI160.XI0.XI0.MM3 N_XI1.XI160.XI0.NET12_XI1.XI160.XI0.XI0.MM3_d
+ N_XI1.G10_XI1.XI160.XI0.XI0.MM3_g
+ N_XI1.XI160.XI0.XI0.NET17_XI1.XI160.XI0.XI0.MM3_s N_VDD_XI1.XI133.XI1.MM3_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=4.125e-13 PD=2.52e-06 PS=5.5e-07
mXI1.XI161.XI0.XI0.MM3 N_XI1.XI161.XI0.NET12_XI1.XI161.XI0.XI0.MM3_d
+ N_XI1.G9_XI1.XI161.XI0.XI0.MM3_g
+ N_XI1.XI161.XI0.XI0.NET17_XI1.XI161.XI0.XI0.MM3_s N_VDD_XI1.XI132.XI1.MM3_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=4.125e-13 PD=2.52e-06 PS=5.5e-07
mXI1.XI162.XI0.XI0.MM3 N_XI1.XI162.XI0.NET12_XI1.XI162.XI0.XI0.MM3_d
+ N_XI1.G8_XI1.XI162.XI0.XI0.MM3_g
+ N_XI1.XI162.XI0.XI0.NET17_XI1.XI162.XI0.XI0.MM3_s N_VDD_XI1.XI131.XI1.MM3_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=4.125e-13 PD=2.52e-06 PS=5.5e-07
mXI1.XI121.XI0.XI0.MM3 N_XI1.XI121.XI0.NET12_XI1.XI121.XI0.XI0.MM3_d
+ N_XI1.G7_XI1.XI121.XI0.XI0.MM3_g
+ N_XI1.XI121.XI0.XI0.NET17_XI1.XI121.XI0.XI0.MM3_s N_VDD_XI1.XI111.XI1.MM3_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=4.125e-13 PD=2.52e-06 PS=5.5e-07
mXI1.XI120.XI0.XI0.MM3 N_XI1.XI120.XI0.NET12_XI1.XI120.XI0.XI0.MM3_d
+ N_XI1.G6_XI1.XI120.XI0.XI0.MM3_g
+ N_XI1.XI120.XI0.XI0.NET17_XI1.XI120.XI0.XI0.MM3_s N_VDD_XI1.XI110.XI1.MM3_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=4.125e-13 PD=2.52e-06 PS=5.5e-07
mXI1.XI119.XI0.XI0.MM3 N_XI1.XI119.XI0.NET12_XI1.XI119.XI0.XI0.MM3_d
+ N_XI1.G5_XI1.XI119.XI0.XI0.MM3_g
+ N_XI1.XI119.XI0.XI0.NET17_XI1.XI119.XI0.XI0.MM3_s N_VDD_XI1.XI103.XI1.MM3_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=4.125e-13 PD=2.52e-06 PS=5.5e-07
mXI1.XI118.XI0.XI0.MM3 N_XI1.XI118.XI0.NET12_XI1.XI118.XI0.XI0.MM3_d
+ N_XI1.G4_XI1.XI118.XI0.XI0.MM3_g
+ N_XI1.XI118.XI0.XI0.NET17_XI1.XI118.XI0.XI0.MM3_s N_VDD_XI1.XI102.XI1.MM3_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=4.125e-13 PD=2.52e-06 PS=5.5e-07
mXI1.XI91.XI0.XI0.MM3 N_XI1.XI91.XI0.NET12_XI1.XI91.XI0.XI0.MM3_d
+ N_XI1.G3_XI1.XI91.XI0.XI0.MM3_g
+ N_XI1.XI91.XI0.XI0.NET17_XI1.XI91.XI0.XI0.MM3_s N_VDD_XI1.XI88.XI1.MM3_b P_18
+ L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=4.125e-13 PD=2.52e-06 PS=5.5e-07
mXI1.XI90.XI0.XI0.MM3 N_XI1.XI90.XI0.NET12_XI1.XI90.XI0.XI0.MM3_d
+ N_XI1.G2_XI1.XI90.XI0.XI0.MM3_g
+ N_XI1.XI90.XI0.XI0.NET17_XI1.XI90.XI0.XI0.MM3_s N_VDD_XI1.XI82.XI1.MM3_b P_18
+ L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=4.125e-13 PD=2.52e-06 PS=5.5e-07
mXI1.XI89.XI0.XI0.MM3 N_XI1.XI89.XI0.NET12_XI1.XI89.XI0.XI0.MM3_d
+ N_XI1.G1_XI1.XI89.XI0.XI0.MM3_g
+ N_XI1.XI89.XI0.XI0.NET17_XI1.XI89.XI0.XI0.MM3_s N_VDD_XI1.XI10.XI1.MM3_b P_18
+ L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=4.125e-13 PD=2.52e-06 PS=5.5e-07
mXI1.XI168.XI0.XI1.MM1 N_XI1.NET198_XI1.XI168.XI0.XI1.MM1_d
+ N_XI1.XI168.XI0.NET12_XI1.XI168.XI0.XI1.MM1_g N_VDD_XI1.XI168.XI0.XI1.MM1_s
+ N_VDD_XI1.XI153.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI1.XI167.XI0.XI1.MM1 N_XI1.NET288_XI1.XI167.XI0.XI1.MM1_d
+ N_XI1.XI167.XI0.NET12_XI1.XI167.XI0.XI1.MM1_g N_VDD_XI1.XI167.XI0.XI1.MM1_s
+ N_VDD_XI1.XI154.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI1.XI166.XI0.XI1.MM1 N_XI1.NET282_XI1.XI166.XI0.XI1.MM1_d
+ N_XI1.XI166.XI0.NET12_XI1.XI166.XI0.XI1.MM1_g N_VDD_XI1.XI166.XI0.XI1.MM1_s
+ N_VDD_XI1.XI157.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI1.XI165.XI0.XI1.MM1 N_XI1.NET276_XI1.XI165.XI0.XI1.MM1_d
+ N_XI1.XI165.XI0.NET12_XI1.XI165.XI0.XI1.MM1_g N_VDD_XI1.XI165.XI0.XI1.MM1_s
+ N_VDD_XI1.XI156.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI1.XI159.XI0.XI1.MM1 N_XI1.NET270_XI1.XI159.XI0.XI1.MM1_d
+ N_XI1.XI159.XI0.NET12_XI1.XI159.XI0.XI1.MM1_g N_VDD_XI1.XI159.XI0.XI1.MM1_s
+ N_VDD_XI1.XI155.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI1.XI160.XI0.XI1.MM1 N_XI1.NET246_XI1.XI160.XI0.XI1.MM1_d
+ N_XI1.XI160.XI0.NET12_XI1.XI160.XI0.XI1.MM1_g N_VDD_XI1.XI160.XI0.XI1.MM1_s
+ N_VDD_XI1.XI133.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI1.XI161.XI0.XI1.MM1 N_XI1.NET252_XI1.XI161.XI0.XI1.MM1_d
+ N_XI1.XI161.XI0.NET12_XI1.XI161.XI0.XI1.MM1_g N_VDD_XI1.XI161.XI0.XI1.MM1_s
+ N_VDD_XI1.XI132.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI1.XI162.XI0.XI1.MM1 N_XI1.NET258_XI1.XI162.XI0.XI1.MM1_d
+ N_XI1.XI162.XI0.NET12_XI1.XI162.XI0.XI1.MM1_g N_VDD_XI1.XI162.XI0.XI1.MM1_s
+ N_VDD_XI1.XI131.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI1.XI121.XI0.XI1.MM1 N_XI1.NET264_XI1.XI121.XI0.XI1.MM1_d
+ N_XI1.XI121.XI0.NET12_XI1.XI121.XI0.XI1.MM1_g N_VDD_XI1.XI121.XI0.XI1.MM1_s
+ N_VDD_XI1.XI111.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI1.XI120.XI0.XI1.MM1 N_XI1.NET204_XI1.XI120.XI0.XI1.MM1_d
+ N_XI1.XI120.XI0.NET12_XI1.XI120.XI0.XI1.MM1_g N_VDD_XI1.XI120.XI0.XI1.MM1_s
+ N_VDD_XI1.XI110.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI1.XI119.XI0.XI1.MM1 N_XI1.NET210_XI1.XI119.XI0.XI1.MM1_d
+ N_XI1.XI119.XI0.NET12_XI1.XI119.XI0.XI1.MM1_g N_VDD_XI1.XI119.XI0.XI1.MM1_s
+ N_VDD_XI1.XI103.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI1.XI118.XI0.XI1.MM1 N_XI1.NET216_XI1.XI118.XI0.XI1.MM1_d
+ N_XI1.XI118.XI0.NET12_XI1.XI118.XI0.XI1.MM1_g N_VDD_XI1.XI118.XI0.XI1.MM1_s
+ N_VDD_XI1.XI102.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI1.XI91.XI0.XI1.MM1 N_XI1.NET222_XI1.XI91.XI0.XI1.MM1_d
+ N_XI1.XI91.XI0.NET12_XI1.XI91.XI0.XI1.MM1_g N_VDD_XI1.XI91.XI0.XI1.MM1_s
+ N_VDD_XI1.XI88.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI1.XI90.XI0.XI1.MM1 N_XI1.NET228_XI1.XI90.XI0.XI1.MM1_d
+ N_XI1.XI90.XI0.NET12_XI1.XI90.XI0.XI1.MM1_g N_VDD_XI1.XI90.XI0.XI1.MM1_s
+ N_VDD_XI1.XI82.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI1.XI89.XI0.XI1.MM1 N_XI1.NET240_XI1.XI89.XI0.XI1.MM1_d
+ N_XI1.XI89.XI0.NET12_XI1.XI89.XI0.XI1.MM1_g N_VDD_XI1.XI89.XI0.XI1.MM1_s
+ N_VDD_XI1.XI10.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13
+ PD=2.48e-06 PS=2.48e-06
mXI19.XI18.MM5 N_XI19.XI18.NET7_XI19.XI18.MM5_d N_NET01249_XI19.XI18.MM5_g
+ N_VDD_XI19.XI18.MM5_s N_VDD_XI1.XI134.XI9.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI19.XI19.MM5 N_XI19.XI19.NET7_XI19.XI19.MM5_d N_NET01249_XI19.XI19.MM5_g
+ N_VDD_XI19.XI19.MM5_s N_VDD_XI1.XI153.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI19.XI17.MM5 N_XI19.XI17.NET7_XI19.XI17.MM5_d N_NET01249_XI19.XI17.MM5_g
+ N_VDD_XI19.XI17.MM5_s N_VDD_XI1.XI154.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI19.XI16.MM5 N_XI19.XI16.NET7_XI19.XI16.MM5_d N_NET01249_XI19.XI16.MM5_g
+ N_VDD_XI19.XI16.MM5_s N_VDD_XI1.XI157.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI19.XI21.MM5 N_XI19.XI21.NET7_XI19.XI21.MM5_d N_NET01249_XI19.XI21.MM5_g
+ N_VDD_XI19.XI21.MM5_s N_VDD_XI1.XI156.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI19.XI20.MM5 N_XI19.XI20.NET7_XI19.XI20.MM5_d N_NET01249_XI19.XI20.MM5_g
+ N_VDD_XI19.XI20.MM5_s N_VDD_XI1.XI155.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI19.XI22.MM5 N_XI19.XI22.NET7_XI19.XI22.MM5_d N_NET01249_XI19.XI22.MM5_g
+ N_VDD_XI19.XI22.MM5_s N_VDD_XI1.XI133.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI19.XI6.MM5 N_XI19.XI6.NET7_XI19.XI6.MM5_d N_NET01249_XI19.XI6.MM5_g
+ N_VDD_XI19.XI6.MM5_s N_VDD_XI1.XI132.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI19.XI5.MM5 N_XI19.XI5.NET7_XI19.XI5.MM5_d N_NET01249_XI19.XI5.MM5_g
+ N_VDD_XI19.XI5.MM5_s N_VDD_XI1.XI131.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI19.XI7.MM5 N_XI19.XI7.NET7_XI19.XI7.MM5_d N_NET01249_XI19.XI7.MM5_g
+ N_VDD_XI19.XI7.MM5_s N_VDD_XI1.XI111.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI19.XI8.MM5 N_XI19.XI8.NET7_XI19.XI8.MM5_d N_NET01249_XI19.XI8.MM5_g
+ N_VDD_XI19.XI8.MM5_s N_VDD_XI1.XI110.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI19.XI3.MM5 N_XI19.XI3.NET7_XI19.XI3.MM5_d N_NET01249_XI19.XI3.MM5_g
+ N_VDD_XI19.XI3.MM5_s N_VDD_XI1.XI103.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI19.XI4.MM5 N_XI19.XI4.NET7_XI19.XI4.MM5_d N_NET01249_XI19.XI4.MM5_g
+ N_VDD_XI19.XI4.MM5_s N_VDD_XI1.XI102.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI19.XI2.MM5 N_XI19.XI2.NET7_XI19.XI2.MM5_d N_NET01249_XI19.XI2.MM5_g
+ N_VDD_XI19.XI2.MM5_s N_VDD_XI1.XI88.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI19.XI1.MM5 N_XI19.XI1.NET7_XI19.XI1.MM5_d N_NET01249_XI19.XI1.MM5_g
+ N_VDD_XI19.XI1.MM5_s N_VDD_XI1.XI82.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI19.XI0.MM5 N_XI19.XI0.NET7_XI19.XI0.MM5_d N_NET01249_XI19.XI0.MM5_g
+ N_VDD_XI19.XI0.MM5_s N_VDD_XI1.XI10.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI19.XI18.MM0 N_NET241_XI19.XI18.MM0_d N_XI19.XI18.NET7_XI19.XI18.MM0_g
+ N_NET559_XI19.XI18.MM0_s N_VDD_XI1.XI134.XI9.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=1.815e-12 AS=9.225e-13 PD=3.92e-06 PS=1.23e-06
mXI19.XI19.MM0 N_NET242_XI19.XI19.MM0_d N_XI19.XI19.NET7_XI19.XI19.MM0_g
+ N_NET560_XI19.XI19.MM0_s N_VDD_XI1.XI153.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=1.815e-12 AS=9.225e-13 PD=3.92e-06 PS=1.23e-06
mXI19.XI17.MM0 N_NET243_XI19.XI17.MM0_d N_XI19.XI17.NET7_XI19.XI17.MM0_g
+ N_NET561_XI19.XI17.MM0_s N_VDD_XI1.XI154.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=1.815e-12 AS=9.225e-13 PD=3.92e-06 PS=1.23e-06
mXI19.XI16.MM0 N_NET244_XI19.XI16.MM0_d N_XI19.XI16.NET7_XI19.XI16.MM0_g
+ N_NET562_XI19.XI16.MM0_s N_VDD_XI1.XI157.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=1.815e-12 AS=9.225e-13 PD=3.92e-06 PS=1.23e-06
mXI19.XI21.MM0 N_NET245_XI19.XI21.MM0_d N_XI19.XI21.NET7_XI19.XI21.MM0_g
+ N_NET563_XI19.XI21.MM0_s N_VDD_XI1.XI156.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=1.815e-12 AS=9.225e-13 PD=3.92e-06 PS=1.23e-06
mXI19.XI20.MM0 N_NET246_XI19.XI20.MM0_d N_XI19.XI20.NET7_XI19.XI20.MM0_g
+ N_NET564_XI19.XI20.MM0_s N_VDD_XI1.XI155.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=1.815e-12 AS=9.225e-13 PD=3.92e-06 PS=1.23e-06
mXI19.XI22.MM0 N_NET247_XI19.XI22.MM0_d N_XI19.XI22.NET7_XI19.XI22.MM0_g
+ N_NET565_XI19.XI22.MM0_s N_VDD_XI1.XI133.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=1.815e-12 AS=9.225e-13 PD=3.92e-06 PS=1.23e-06
mXI19.XI6.MM0 N_NET248_XI19.XI6.MM0_d N_XI19.XI6.NET7_XI19.XI6.MM0_g
+ N_NET566_XI19.XI6.MM0_s N_VDD_XI1.XI132.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=1.815e-12 AS=9.225e-13 PD=3.92e-06 PS=1.23e-06
mXI19.XI5.MM0 N_NET249_XI19.XI5.MM0_d N_XI19.XI5.NET7_XI19.XI5.MM0_g
+ N_NET567_XI19.XI5.MM0_s N_VDD_XI1.XI131.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=1.815e-12 AS=9.225e-13 PD=3.92e-06 PS=1.23e-06
mXI19.XI7.MM0 N_NET250_XI19.XI7.MM0_d N_XI19.XI7.NET7_XI19.XI7.MM0_g
+ N_NET568_XI19.XI7.MM0_s N_VDD_XI1.XI111.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=1.815e-12 AS=9.225e-13 PD=3.92e-06 PS=1.23e-06
mXI19.XI8.MM0 N_NET251_XI19.XI8.MM0_d N_XI19.XI8.NET7_XI19.XI8.MM0_g
+ N_NET569_XI19.XI8.MM0_s N_VDD_XI1.XI110.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=1.815e-12 AS=9.225e-13 PD=3.92e-06 PS=1.23e-06
mXI19.XI3.MM0 N_NET252_XI19.XI3.MM0_d N_XI19.XI3.NET7_XI19.XI3.MM0_g
+ N_NET570_XI19.XI3.MM0_s N_VDD_XI1.XI103.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=1.815e-12 AS=9.225e-13 PD=3.92e-06 PS=1.23e-06
mXI19.XI4.MM0 N_NET253_XI19.XI4.MM0_d N_XI19.XI4.NET7_XI19.XI4.MM0_g
+ N_NET571_XI19.XI4.MM0_s N_VDD_XI1.XI102.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=1.815e-12 AS=9.225e-13 PD=3.92e-06 PS=1.23e-06
mXI19.XI2.MM0 N_NET254_XI19.XI2.MM0_d N_XI19.XI2.NET7_XI19.XI2.MM0_g
+ N_NET572_XI19.XI2.MM0_s N_VDD_XI1.XI88.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=1.815e-12 AS=9.225e-13 PD=3.92e-06 PS=1.23e-06
mXI19.XI1.MM0 N_NET255_XI19.XI1.MM0_d N_XI19.XI1.NET7_XI19.XI1.MM0_g
+ N_NET573_XI19.XI1.MM0_s N_VDD_XI1.XI82.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=1.815e-12 AS=9.225e-13 PD=3.92e-06 PS=1.23e-06
mXI19.XI0.MM0 N_NET256_XI19.XI0.MM0_d N_XI19.XI0.NET7_XI19.XI0.MM0_g
+ N_NET574_XI19.XI0.MM0_s N_VDD_XI1.XI10.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=1.815e-12 AS=9.225e-13 PD=3.92e-06 PS=1.23e-06
mXI19.XI18.MM1 N_MAX15_XI19.XI18.MM1_d N_NET01249_XI19.XI18.MM1_g
+ N_NET559_XI19.XI18.MM1_s N_VDD_XI1.XI134.XI9.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=9.225e-13 PD=2.48e-06 PS=1.23e-06
mXI19.XI19.MM1 N_MAX14_XI19.XI19.MM1_d N_NET01249_XI19.XI19.MM1_g
+ N_NET560_XI19.XI19.MM1_s N_VDD_XI1.XI153.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=9.225e-13 PD=2.48e-06 PS=1.23e-06
mXI19.XI17.MM1 N_MAX13_XI19.XI17.MM1_d N_NET01249_XI19.XI17.MM1_g
+ N_NET561_XI19.XI17.MM1_s N_VDD_XI1.XI154.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=9.225e-13 PD=2.48e-06 PS=1.23e-06
mXI19.XI16.MM1 N_MAX12_XI19.XI16.MM1_d N_NET01249_XI19.XI16.MM1_g
+ N_NET562_XI19.XI16.MM1_s N_VDD_XI1.XI157.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=9.225e-13 PD=2.48e-06 PS=1.23e-06
mXI19.XI21.MM1 N_MAX11_XI19.XI21.MM1_d N_NET01249_XI19.XI21.MM1_g
+ N_NET563_XI19.XI21.MM1_s N_VDD_XI1.XI156.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=9.225e-13 PD=2.48e-06 PS=1.23e-06
mXI19.XI20.MM1 N_MAX10_XI19.XI20.MM1_d N_NET01249_XI19.XI20.MM1_g
+ N_NET564_XI19.XI20.MM1_s N_VDD_XI1.XI155.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=9.225e-13 PD=2.48e-06 PS=1.23e-06
mXI19.XI22.MM1 N_MAX9_XI19.XI22.MM1_d N_NET01249_XI19.XI22.MM1_g
+ N_NET565_XI19.XI22.MM1_s N_VDD_XI1.XI133.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=9.225e-13 PD=2.48e-06 PS=1.23e-06
mXI19.XI6.MM1 N_MAX8_XI19.XI6.MM1_d N_NET01249_XI19.XI6.MM1_g
+ N_NET566_XI19.XI6.MM1_s N_VDD_XI1.XI132.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=9.225e-13 PD=2.48e-06 PS=1.23e-06
mXI19.XI5.MM1 N_MAX7_XI19.XI5.MM1_d N_NET01249_XI19.XI5.MM1_g
+ N_NET567_XI19.XI5.MM1_s N_VDD_XI1.XI131.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=9.225e-13 PD=2.48e-06 PS=1.23e-06
mXI19.XI7.MM1 N_MAX6_XI19.XI7.MM1_d N_NET01249_XI19.XI7.MM1_g
+ N_NET568_XI19.XI7.MM1_s N_VDD_XI1.XI111.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=9.225e-13 PD=2.48e-06 PS=1.23e-06
mXI19.XI8.MM1 N_MAX5_XI19.XI8.MM1_d N_NET01249_XI19.XI8.MM1_g
+ N_NET569_XI19.XI8.MM1_s N_VDD_XI1.XI110.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=9.225e-13 PD=2.48e-06 PS=1.23e-06
mXI19.XI3.MM1 N_MAX4_XI19.XI3.MM1_d N_NET01249_XI19.XI3.MM1_g
+ N_NET570_XI19.XI3.MM1_s N_VDD_XI1.XI103.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=9.225e-13 PD=2.48e-06 PS=1.23e-06
mXI19.XI4.MM1 N_MAX3_XI19.XI4.MM1_d N_NET01249_XI19.XI4.MM1_g
+ N_NET571_XI19.XI4.MM1_s N_VDD_XI1.XI102.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=9.225e-13 PD=2.48e-06 PS=1.23e-06
mXI19.XI2.MM1 N_MAX2_XI19.XI2.MM1_d N_NET01249_XI19.XI2.MM1_g
+ N_NET572_XI19.XI2.MM1_s N_VDD_XI1.XI88.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=9.225e-13 PD=2.48e-06 PS=1.23e-06
mXI19.XI1.MM1 N_MAX1_XI19.XI1.MM1_d N_NET01249_XI19.XI1.MM1_g
+ N_NET573_XI19.XI1.MM1_s N_VDD_XI1.XI82.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=9.225e-13 PD=2.48e-06 PS=1.23e-06
mXI19.XI0.MM1 N_MAX0_XI19.XI0.MM1_d N_NET01249_XI19.XI0.MM1_g
+ N_NET574_XI19.XI0.MM1_s N_VDD_XI1.XI10.XI1.MM3_b P_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=9.225e-13 PD=2.48e-06 PS=1.23e-06
mXI14.MM0 N_XI14.NET116_XI14.MM0_d N_NET198_XI14.MM0_g N_VDD_XI14.MM0_s
+ N_VDD_XI14.MM0_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06
+ PS=2.48e-06
mXI14.XI16.XI0.MM3 N_XI14.XI16.XI0.NET17_XI14.XI16.XI0.MM3_d
+ N_XI14.NET116_XI14.XI16.XI0.MM3_g N_VDD_XI14.XI16.XI0.MM3_s N_VDD_XI14.MM0_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=5.625e-13 AS=7.35e-13 PD=7.5e-07 PS=2.48e-06
mXI14.XI16.XI0.MM1 N_XI14.XI16.NET12_XI14.XI16.XI0.MM1_d
+ N_NET559_XI14.XI16.XI0.MM1_g N_XI14.XI16.XI0.NET17_XI14.XI16.XI0.MM1_s
+ N_VDD_XI14.MM0_b P_18 L=1.8e-07 W=1.5e-06 AD=7.65e-13 AS=5.625e-13 PD=2.52e-06
+ PS=7.5e-07
mXI14.XI16.XI1.MM1 N_NET382_XI14.XI16.XI1.MM1_d
+ N_XI14.XI16.NET12_XI14.XI16.XI1.MM1_g N_VDD_XI14.XI16.XI1.MM1_s
+ N_VDD_XI14.MM0_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06
+ PS=2.48e-06
mXI14.XI15.XI1.MM3 N_XI14.XI15.NET6_XI14.XI15.XI1.MM3_d
+ N_NET198_XI14.XI15.XI1.MM3_g N_VDD_XI14.XI15.XI1.MM3_s N_VDD_XI14.MM0_b P_18
+ L=1.8e-07 W=1.5e-06 AD=4.125e-13 AS=7.35e-13 PD=5.5e-07 PS=2.48e-06
mXI14.XI15.XI1.MM1 N_XI14.XI15.NET6_XI14.XI15.XI1.MM1_d
+ N_NET560_XI14.XI15.XI1.MM1_g N_VDD_XI14.XI15.XI1.MM1_s N_VDD_XI14.MM0_b P_18
+ L=1.8e-07 W=1.5e-06 AD=4.125e-13 AS=7.65e-13 PD=5.5e-07 PS=2.52e-06
mXI14.XI15.XI0.MM1 N_NET383_XI14.XI15.XI0.MM1_d
+ N_XI14.XI15.NET6_XI14.XI15.XI0.MM1_g N_VDD_XI14.XI15.XI0.MM1_s
+ N_VDD_XI14.MM0_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06
+ PS=2.48e-06
mXI14.XI14.XI1.MM3 N_XI14.XI14.NET6_XI14.XI14.XI1.MM3_d
+ N_NET198_XI14.XI14.XI1.MM3_g N_VDD_XI14.XI14.XI1.MM3_s N_VDD_XI14.MM0_b P_18
+ L=1.8e-07 W=1.5e-06 AD=4.125e-13 AS=7.35e-13 PD=5.5e-07 PS=2.48e-06
mXI14.XI14.XI1.MM1 N_XI14.XI14.NET6_XI14.XI14.XI1.MM1_d
+ N_NET561_XI14.XI14.XI1.MM1_g N_VDD_XI14.XI14.XI1.MM1_s N_VDD_XI14.MM0_b P_18
+ L=1.8e-07 W=1.5e-06 AD=4.125e-13 AS=7.65e-13 PD=5.5e-07 PS=2.52e-06
mXI14.XI14.XI0.MM1 N_NET384_XI14.XI14.XI0.MM1_d
+ N_XI14.XI14.NET6_XI14.XI14.XI0.MM1_g N_VDD_XI14.XI14.XI0.MM1_s
+ N_VDD_XI14.MM0_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06
+ PS=2.48e-06
mXI14.XI13.XI1.MM3 N_XI14.XI13.NET6_XI14.XI13.XI1.MM3_d
+ N_NET198_XI14.XI13.XI1.MM3_g N_VDD_XI14.XI13.XI1.MM3_s N_VDD_XI14.MM0_b P_18
+ L=1.8e-07 W=1.5e-06 AD=4.125e-13 AS=7.35e-13 PD=5.5e-07 PS=2.48e-06
mXI14.XI13.XI1.MM1 N_XI14.XI13.NET6_XI14.XI13.XI1.MM1_d
+ N_NET562_XI14.XI13.XI1.MM1_g N_VDD_XI14.XI13.XI1.MM1_s N_VDD_XI14.MM0_b P_18
+ L=1.8e-07 W=1.5e-06 AD=4.125e-13 AS=7.65e-13 PD=5.5e-07 PS=2.52e-06
mXI14.XI13.XI0.MM1 N_NET385_XI14.XI13.XI0.MM1_d
+ N_XI14.XI13.NET6_XI14.XI13.XI0.MM1_g N_VDD_XI14.XI13.XI0.MM1_s
+ N_VDD_XI14.MM0_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06
+ PS=2.48e-06
mXI14.XI12.XI1.MM3 N_XI14.XI12.NET6_XI14.XI12.XI1.MM3_d
+ N_NET198_XI14.XI12.XI1.MM3_g N_VDD_XI14.XI12.XI1.MM3_s N_VDD_XI14.MM0_b P_18
+ L=1.8e-07 W=1.5e-06 AD=4.125e-13 AS=7.35e-13 PD=5.5e-07 PS=2.48e-06
mXI14.XI12.XI1.MM1 N_XI14.XI12.NET6_XI14.XI12.XI1.MM1_d
+ N_NET563_XI14.XI12.XI1.MM1_g N_VDD_XI14.XI12.XI1.MM1_s N_VDD_XI14.MM0_b P_18
+ L=1.8e-07 W=1.5e-06 AD=4.125e-13 AS=7.65e-13 PD=5.5e-07 PS=2.52e-06
mXI14.XI12.XI0.MM1 N_NET386_XI14.XI12.XI0.MM1_d
+ N_XI14.XI12.NET6_XI14.XI12.XI0.MM1_g N_VDD_XI14.XI12.XI0.MM1_s
+ N_VDD_XI14.MM0_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06
+ PS=2.48e-06
mXI14.XI11.XI1.MM3 N_XI14.XI11.NET6_XI14.XI11.XI1.MM3_d
+ N_NET198_XI14.XI11.XI1.MM3_g N_VDD_XI14.XI11.XI1.MM3_s N_VDD_XI14.MM0_b P_18
+ L=1.8e-07 W=1.5e-06 AD=4.125e-13 AS=7.35e-13 PD=5.5e-07 PS=2.48e-06
mXI14.XI11.XI1.MM1 N_XI14.XI11.NET6_XI14.XI11.XI1.MM1_d
+ N_NET564_XI14.XI11.XI1.MM1_g N_VDD_XI14.XI11.XI1.MM1_s N_VDD_XI14.MM0_b P_18
+ L=1.8e-07 W=1.5e-06 AD=4.125e-13 AS=7.65e-13 PD=5.5e-07 PS=2.52e-06
mXI14.XI11.XI0.MM1 N_NET387_XI14.XI11.XI0.MM1_d
+ N_XI14.XI11.NET6_XI14.XI11.XI0.MM1_g N_VDD_XI14.XI11.XI0.MM1_s
+ N_VDD_XI14.MM0_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06
+ PS=2.48e-06
mXI14.XI10.XI1.MM3 N_XI14.XI10.NET6_XI14.XI10.XI1.MM3_d
+ N_NET198_XI14.XI10.XI1.MM3_g N_VDD_XI14.XI10.XI1.MM3_s N_VDD_XI14.MM0_b P_18
+ L=1.8e-07 W=1.5e-06 AD=4.125e-13 AS=7.35e-13 PD=5.5e-07 PS=2.48e-06
mXI14.XI10.XI1.MM1 N_XI14.XI10.NET6_XI14.XI10.XI1.MM1_d
+ N_NET565_XI14.XI10.XI1.MM1_g N_VDD_XI14.XI10.XI1.MM1_s N_VDD_XI14.MM0_b P_18
+ L=1.8e-07 W=1.5e-06 AD=4.125e-13 AS=7.65e-13 PD=5.5e-07 PS=2.52e-06
mXI14.XI10.XI0.MM1 N_NET388_XI14.XI10.XI0.MM1_d
+ N_XI14.XI10.NET6_XI14.XI10.XI0.MM1_g N_VDD_XI14.XI10.XI0.MM1_s
+ N_VDD_XI14.MM0_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=7.35e-13 PD=2.48e-06
+ PS=2.48e-06
mXI14.XI9.XI1.MM3 N_XI14.XI9.NET6_XI14.XI9.XI1.MM3_d N_NET198_XI14.XI9.XI1.MM3_g
+ N_VDD_XI14.XI9.XI1.MM3_s N_VDD_XI14.MM0_b P_18 L=1.8e-07 W=1.5e-06
+ AD=4.125e-13 AS=7.35e-13 PD=5.5e-07 PS=2.48e-06
mXI14.XI9.XI1.MM1 N_XI14.XI9.NET6_XI14.XI9.XI1.MM1_d N_NET566_XI14.XI9.XI1.MM1_g
+ N_VDD_XI14.XI9.XI1.MM1_s N_VDD_XI14.MM0_b P_18 L=1.8e-07 W=1.5e-06
+ AD=4.125e-13 AS=7.65e-13 PD=5.5e-07 PS=2.52e-06
mXI14.XI9.XI0.MM1 N_NET389_XI14.XI9.XI0.MM1_d N_XI14.XI9.NET6_XI14.XI9.XI0.MM1_g
+ N_VDD_XI14.XI9.XI0.MM1_s N_VDD_XI14.MM0_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13
+ AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI14.XI8.XI1.MM3 N_XI14.XI8.NET6_XI14.XI8.XI1.MM3_d N_NET198_XI14.XI8.XI1.MM3_g
+ N_VDD_XI14.XI8.XI1.MM3_s N_VDD_XI14.MM0_b P_18 L=1.8e-07 W=1.5e-06
+ AD=4.125e-13 AS=7.35e-13 PD=5.5e-07 PS=2.48e-06
mXI14.XI8.XI1.MM1 N_XI14.XI8.NET6_XI14.XI8.XI1.MM1_d N_NET567_XI14.XI8.XI1.MM1_g
+ N_VDD_XI14.XI8.XI1.MM1_s N_VDD_XI14.MM0_b P_18 L=1.8e-07 W=1.5e-06
+ AD=4.125e-13 AS=7.65e-13 PD=5.5e-07 PS=2.52e-06
mXI14.XI8.XI0.MM1 N_NET390_XI14.XI8.XI0.MM1_d N_XI14.XI8.NET6_XI14.XI8.XI0.MM1_g
+ N_VDD_XI14.XI8.XI0.MM1_s N_VDD_XI14.MM0_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13
+ AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI14.XI7.XI1.MM3 N_XI14.XI7.NET6_XI14.XI7.XI1.MM3_d N_NET198_XI14.XI7.XI1.MM3_g
+ N_VDD_XI14.XI7.XI1.MM3_s N_VDD_XI14.MM0_b P_18 L=1.8e-07 W=1.5e-06
+ AD=4.125e-13 AS=7.35e-13 PD=5.5e-07 PS=2.48e-06
mXI14.XI7.XI1.MM1 N_XI14.XI7.NET6_XI14.XI7.XI1.MM1_d N_NET568_XI14.XI7.XI1.MM1_g
+ N_VDD_XI14.XI7.XI1.MM1_s N_VDD_XI14.MM0_b P_18 L=1.8e-07 W=1.5e-06
+ AD=4.125e-13 AS=7.65e-13 PD=5.5e-07 PS=2.52e-06
mXI14.XI7.XI0.MM1 N_NET391_XI14.XI7.XI0.MM1_d N_XI14.XI7.NET6_XI14.XI7.XI0.MM1_g
+ N_VDD_XI14.XI7.XI0.MM1_s N_VDD_XI14.MM0_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13
+ AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI14.XI6.XI1.MM3 N_XI14.XI6.NET6_XI14.XI6.XI1.MM3_d N_NET198_XI14.XI6.XI1.MM3_g
+ N_VDD_XI14.XI6.XI1.MM3_s N_VDD_XI14.MM0_b P_18 L=1.8e-07 W=1.5e-06
+ AD=4.125e-13 AS=7.35e-13 PD=5.5e-07 PS=2.48e-06
mXI14.XI6.XI1.MM1 N_XI14.XI6.NET6_XI14.XI6.XI1.MM1_d N_NET569_XI14.XI6.XI1.MM1_g
+ N_VDD_XI14.XI6.XI1.MM1_s N_VDD_XI14.MM0_b P_18 L=1.8e-07 W=1.5e-06
+ AD=4.125e-13 AS=7.65e-13 PD=5.5e-07 PS=2.52e-06
mXI14.XI6.XI0.MM1 N_NET392_XI14.XI6.XI0.MM1_d N_XI14.XI6.NET6_XI14.XI6.XI0.MM1_g
+ N_VDD_XI14.XI6.XI0.MM1_s N_VDD_XI14.MM0_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13
+ AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI14.XI5.XI1.MM3 N_XI14.XI5.NET6_XI14.XI5.XI1.MM3_d N_NET198_XI14.XI5.XI1.MM3_g
+ N_VDD_XI14.XI5.XI1.MM3_s N_VDD_XI14.MM0_b P_18 L=1.8e-07 W=1.5e-06
+ AD=4.125e-13 AS=7.35e-13 PD=5.5e-07 PS=2.48e-06
mXI14.XI5.XI1.MM1 N_XI14.XI5.NET6_XI14.XI5.XI1.MM1_d N_NET570_XI14.XI5.XI1.MM1_g
+ N_VDD_XI14.XI5.XI1.MM1_s N_VDD_XI14.MM0_b P_18 L=1.8e-07 W=1.5e-06
+ AD=4.125e-13 AS=7.65e-13 PD=5.5e-07 PS=2.52e-06
mXI14.XI5.XI0.MM1 N_NET393_XI14.XI5.XI0.MM1_d N_XI14.XI5.NET6_XI14.XI5.XI0.MM1_g
+ N_VDD_XI14.XI5.XI0.MM1_s N_VDD_XI14.MM0_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13
+ AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI14.XI4.XI1.MM3 N_XI14.XI4.NET6_XI14.XI4.XI1.MM3_d N_NET198_XI14.XI4.XI1.MM3_g
+ N_VDD_XI14.XI4.XI1.MM3_s N_VDD_XI14.MM0_b P_18 L=1.8e-07 W=1.5e-06
+ AD=4.125e-13 AS=7.35e-13 PD=5.5e-07 PS=2.48e-06
mXI14.XI4.XI1.MM1 N_XI14.XI4.NET6_XI14.XI4.XI1.MM1_d N_NET571_XI14.XI4.XI1.MM1_g
+ N_VDD_XI14.XI4.XI1.MM1_s N_VDD_XI14.MM0_b P_18 L=1.8e-07 W=1.5e-06
+ AD=4.125e-13 AS=7.65e-13 PD=5.5e-07 PS=2.52e-06
mXI14.XI4.XI0.MM1 N_NET394_XI14.XI4.XI0.MM1_d N_XI14.XI4.NET6_XI14.XI4.XI0.MM1_g
+ N_VDD_XI14.XI4.XI0.MM1_s N_VDD_XI14.MM0_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13
+ AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI14.XI3.XI1.MM3 N_XI14.XI3.NET6_XI14.XI3.XI1.MM3_d N_NET198_XI14.XI3.XI1.MM3_g
+ N_VDD_XI14.XI3.XI1.MM3_s N_VDD_XI14.MM0_b P_18 L=1.8e-07 W=1.5e-06
+ AD=4.125e-13 AS=7.35e-13 PD=5.5e-07 PS=2.48e-06
mXI14.XI3.XI1.MM1 N_XI14.XI3.NET6_XI14.XI3.XI1.MM1_d N_NET572_XI14.XI3.XI1.MM1_g
+ N_VDD_XI14.XI3.XI1.MM1_s N_VDD_XI14.MM0_b P_18 L=1.8e-07 W=1.5e-06
+ AD=4.125e-13 AS=7.65e-13 PD=5.5e-07 PS=2.52e-06
mXI14.XI3.XI0.MM1 N_NET395_XI14.XI3.XI0.MM1_d N_XI14.XI3.NET6_XI14.XI3.XI0.MM1_g
+ N_VDD_XI14.XI3.XI0.MM1_s N_VDD_XI14.MM0_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13
+ AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI14.XI2.XI1.MM3 N_XI14.XI2.NET6_XI14.XI2.XI1.MM3_d N_NET198_XI14.XI2.XI1.MM3_g
+ N_VDD_XI14.XI2.XI1.MM3_s N_VDD_XI14.MM0_b P_18 L=1.8e-07 W=1.5e-06
+ AD=4.125e-13 AS=7.35e-13 PD=5.5e-07 PS=2.48e-06
mXI14.XI2.XI1.MM1 N_XI14.XI2.NET6_XI14.XI2.XI1.MM1_d N_NET573_XI14.XI2.XI1.MM1_g
+ N_VDD_XI14.XI2.XI1.MM1_s N_VDD_XI14.MM0_b P_18 L=1.8e-07 W=1.5e-06
+ AD=4.125e-13 AS=7.65e-13 PD=5.5e-07 PS=2.52e-06
mXI14.XI2.XI0.MM1 N_NET396_XI14.XI2.XI0.MM1_d N_XI14.XI2.NET6_XI14.XI2.XI0.MM1_g
+ N_VDD_XI14.XI2.XI0.MM1_s N_VDD_XI14.MM0_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13
+ AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI14.XI1.XI1.MM3 N_XI14.XI1.NET6_XI14.XI1.XI1.MM3_d N_NET198_XI14.XI1.XI1.MM3_g
+ N_VDD_XI14.XI1.XI1.MM3_s N_VDD_XI14.MM0_b P_18 L=1.8e-07 W=1.5e-06
+ AD=4.125e-13 AS=7.35e-13 PD=5.5e-07 PS=2.48e-06
mXI14.XI1.XI1.MM1 N_XI14.XI1.NET6_XI14.XI1.XI1.MM1_d N_NET574_XI14.XI1.XI1.MM1_g
+ N_VDD_XI14.XI1.XI1.MM1_s N_VDD_XI14.MM0_b P_18 L=1.8e-07 W=1.5e-06
+ AD=4.125e-13 AS=7.65e-13 PD=5.5e-07 PS=2.52e-06
mXI14.XI1.XI0.MM1 N_NET397_XI14.XI1.XI0.MM1_d N_XI14.XI1.NET6_XI14.XI1.XI0.MM1_g
+ N_VDD_XI14.XI1.XI0.MM1_s N_VDD_XI14.MM0_b P_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13
+ AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI13.XI30.XI0.MM1 N_XI13.XI30.NET0180_XI13.XI30.XI0.MM1_d
+ N_NET222_XI13.XI30.XI0.MM1_g N_VDD_XI13.XI30.XI0.MM1_s
+ N_VDD_XI13.XI30.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI13.XI29.XI0.MM1 N_XI13.XI29.NET0180_XI13.XI29.XI0.MM1_d
+ N_NET222_XI13.XI29.XI0.MM1_g N_VDD_XI13.XI29.XI0.MM1_s
+ N_VDD_XI13.XI29.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI13.XI31.XI0.MM1 N_XI13.XI31.NET0180_XI13.XI31.XI0.MM1_d
+ N_NET222_XI13.XI31.XI0.MM1_g N_VDD_XI13.XI31.XI0.MM1_s
+ N_VDD_XI13.XI31.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI13.XI28.XI0.MM1 N_XI13.XI28.NET0180_XI13.XI28.XI0.MM1_d
+ N_NET222_XI13.XI28.XI0.MM1_g N_VDD_XI13.XI28.XI0.MM1_s
+ N_VDD_XI13.XI28.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI13.XI25.XI0.MM1 N_XI13.XI25.NET0180_XI13.XI25.XI0.MM1_d
+ N_NET222_XI13.XI25.XI0.MM1_g N_VDD_XI13.XI25.XI0.MM1_s
+ N_VDD_XI13.XI25.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI13.XI26.XI0.MM1 N_XI13.XI26.NET0180_XI13.XI26.XI0.MM1_d
+ N_NET222_XI13.XI26.XI0.MM1_g N_VDD_XI13.XI26.XI0.MM1_s
+ N_VDD_XI13.XI26.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI13.XI24.XI0.MM1 N_XI13.XI24.NET0180_XI13.XI24.XI0.MM1_d
+ N_NET222_XI13.XI24.XI0.MM1_g N_VDD_XI13.XI24.XI0.MM1_s
+ N_VDD_XI13.XI24.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI13.XI27.XI0.MM1 N_XI13.XI27.NET0180_XI13.XI27.XI0.MM1_d
+ N_NET222_XI13.XI27.XI0.MM1_g N_VDD_XI13.XI27.XI0.MM1_s
+ N_VDD_XI13.XI27.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI13.XI22.XI0.MM1 N_XI13.XI22.NET0180_XI13.XI22.XI0.MM1_d
+ N_NET222_XI13.XI22.XI0.MM1_g N_VDD_XI13.XI22.XI0.MM1_s
+ N_VDD_XI13.XI22.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI13.XI21.XI0.MM1 N_XI13.XI21.NET0180_XI13.XI21.XI0.MM1_d
+ N_NET222_XI13.XI21.XI0.MM1_g N_VDD_XI13.XI21.XI0.MM1_s
+ N_VDD_XI13.XI21.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI13.XI23.XI0.MM1 N_XI13.XI23.NET0180_XI13.XI23.XI0.MM1_d
+ N_NET222_XI13.XI23.XI0.MM1_g N_VDD_XI13.XI23.XI0.MM1_s
+ N_VDD_XI13.XI23.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI13.XI19.XI0.MM1 N_XI13.XI19.NET0180_XI13.XI19.XI0.MM1_d
+ N_NET222_XI13.XI19.XI0.MM1_g N_VDD_XI13.XI19.XI0.MM1_s
+ N_VDD_XI13.XI19.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI13.XI20.XI0.MM1 N_XI13.XI20.NET0180_XI13.XI20.XI0.MM1_d
+ N_NET222_XI13.XI20.XI0.MM1_g N_VDD_XI13.XI20.XI0.MM1_s
+ N_VDD_XI13.XI20.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI13.XI18.XI0.MM1 N_XI13.XI18.NET0180_XI13.XI18.XI0.MM1_d
+ N_NET222_XI13.XI18.XI0.MM1_g N_VDD_XI13.XI18.XI0.MM1_s
+ N_VDD_XI13.XI18.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI13.XI17.XI0.MM1 N_XI13.XI17.NET0180_XI13.XI17.XI0.MM1_d
+ N_NET222_XI13.XI17.XI0.MM1_g N_VDD_XI13.XI17.XI0.MM1_s
+ N_VDD_XI13.XI17.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI13.XI0.XI0.MM1 N_XI13.XI0.NET0180_XI13.XI0.XI0.MM1_d
+ N_NET222_XI13.XI0.XI0.MM1_g N_VDD_XI13.XI0.XI0.MM1_s N_VDD_XI13.XI0.XI0.MM1_b
+ P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI13.XI30.XI1.MM1 N_XI13.XI30.NET35_XI13.XI30.XI1.MM1_d
+ N_XI13.XI30.NET0180_XI13.XI30.XI1.MM1_g N_VDD_XI13.XI30.XI1.MM1_s
+ N_VDD_XI13.XI30.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI13.XI29.XI1.MM1 N_XI13.XI29.NET35_XI13.XI29.XI1.MM1_d
+ N_XI13.XI29.NET0180_XI13.XI29.XI1.MM1_g N_VDD_XI13.XI29.XI1.MM1_s
+ N_VDD_XI13.XI29.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI13.XI31.XI1.MM1 N_XI13.XI31.NET35_XI13.XI31.XI1.MM1_d
+ N_XI13.XI31.NET0180_XI13.XI31.XI1.MM1_g N_VDD_XI13.XI31.XI1.MM1_s
+ N_VDD_XI13.XI31.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI13.XI28.XI1.MM1 N_XI13.XI28.NET35_XI13.XI28.XI1.MM1_d
+ N_XI13.XI28.NET0180_XI13.XI28.XI1.MM1_g N_VDD_XI13.XI28.XI1.MM1_s
+ N_VDD_XI13.XI28.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI13.XI25.XI1.MM1 N_XI13.XI25.NET35_XI13.XI25.XI1.MM1_d
+ N_XI13.XI25.NET0180_XI13.XI25.XI1.MM1_g N_VDD_XI13.XI25.XI1.MM1_s
+ N_VDD_XI13.XI25.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI13.XI26.XI1.MM1 N_XI13.XI26.NET35_XI13.XI26.XI1.MM1_d
+ N_XI13.XI26.NET0180_XI13.XI26.XI1.MM1_g N_VDD_XI13.XI26.XI1.MM1_s
+ N_VDD_XI13.XI26.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI13.XI24.XI1.MM1 N_XI13.XI24.NET35_XI13.XI24.XI1.MM1_d
+ N_XI13.XI24.NET0180_XI13.XI24.XI1.MM1_g N_VDD_XI13.XI24.XI1.MM1_s
+ N_VDD_XI13.XI24.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI13.XI27.XI1.MM1 N_XI13.XI27.NET35_XI13.XI27.XI1.MM1_d
+ N_XI13.XI27.NET0180_XI13.XI27.XI1.MM1_g N_VDD_XI13.XI27.XI1.MM1_s
+ N_VDD_XI13.XI27.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI13.XI22.XI1.MM1 N_XI13.XI22.NET35_XI13.XI22.XI1.MM1_d
+ N_XI13.XI22.NET0180_XI13.XI22.XI1.MM1_g N_VDD_XI13.XI22.XI1.MM1_s
+ N_VDD_XI13.XI22.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI13.XI21.XI1.MM1 N_XI13.XI21.NET35_XI13.XI21.XI1.MM1_d
+ N_XI13.XI21.NET0180_XI13.XI21.XI1.MM1_g N_VDD_XI13.XI21.XI1.MM1_s
+ N_VDD_XI13.XI21.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI13.XI23.XI1.MM1 N_XI13.XI23.NET35_XI13.XI23.XI1.MM1_d
+ N_XI13.XI23.NET0180_XI13.XI23.XI1.MM1_g N_VDD_XI13.XI23.XI1.MM1_s
+ N_VDD_XI13.XI23.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI13.XI19.XI1.MM1 N_XI13.XI19.NET35_XI13.XI19.XI1.MM1_d
+ N_XI13.XI19.NET0180_XI13.XI19.XI1.MM1_g N_VDD_XI13.XI19.XI1.MM1_s
+ N_VDD_XI13.XI19.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI13.XI20.XI1.MM1 N_XI13.XI20.NET35_XI13.XI20.XI1.MM1_d
+ N_XI13.XI20.NET0180_XI13.XI20.XI1.MM1_g N_VDD_XI13.XI20.XI1.MM1_s
+ N_VDD_XI13.XI20.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI13.XI18.XI1.MM1 N_XI13.XI18.NET35_XI13.XI18.XI1.MM1_d
+ N_XI13.XI18.NET0180_XI13.XI18.XI1.MM1_g N_VDD_XI13.XI18.XI1.MM1_s
+ N_VDD_XI13.XI18.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI13.XI17.XI1.MM1 N_XI13.XI17.NET35_XI13.XI17.XI1.MM1_d
+ N_XI13.XI17.NET0180_XI13.XI17.XI1.MM1_g N_VDD_XI13.XI17.XI1.MM1_s
+ N_VDD_XI13.XI17.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI13.XI0.XI1.MM1 N_XI13.XI0.NET35_XI13.XI0.XI1.MM1_d
+ N_XI13.XI0.NET0180_XI13.XI0.XI1.MM1_g N_VDD_XI13.XI0.XI1.MM1_s
+ N_VDD_XI13.XI0.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI13.XI30.MM25 N_XI13.XI30.CLKB_XI13.XI30.MM25_d
+ N_XI13.XI30.NET35_XI13.XI30.MM25_g N_VDD_XI13.XI30.MM25_s
+ N_VDD_XI13.XI30.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI13.XI29.MM25 N_XI13.XI29.CLKB_XI13.XI29.MM25_d
+ N_XI13.XI29.NET35_XI13.XI29.MM25_g N_VDD_XI13.XI29.MM25_s
+ N_VDD_XI13.XI29.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI13.XI31.MM25 N_XI13.XI31.CLKB_XI13.XI31.MM25_d
+ N_XI13.XI31.NET35_XI13.XI31.MM25_g N_VDD_XI13.XI31.MM25_s
+ N_VDD_XI13.XI31.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI13.XI28.MM25 N_XI13.XI28.CLKB_XI13.XI28.MM25_d
+ N_XI13.XI28.NET35_XI13.XI28.MM25_g N_VDD_XI13.XI28.MM25_s
+ N_VDD_XI13.XI28.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI13.XI25.MM25 N_XI13.XI25.CLKB_XI13.XI25.MM25_d
+ N_XI13.XI25.NET35_XI13.XI25.MM25_g N_VDD_XI13.XI25.MM25_s
+ N_VDD_XI13.XI25.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI13.XI26.MM25 N_XI13.XI26.CLKB_XI13.XI26.MM25_d
+ N_XI13.XI26.NET35_XI13.XI26.MM25_g N_VDD_XI13.XI26.MM25_s
+ N_VDD_XI13.XI26.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI13.XI24.MM25 N_XI13.XI24.CLKB_XI13.XI24.MM25_d
+ N_XI13.XI24.NET35_XI13.XI24.MM25_g N_VDD_XI13.XI24.MM25_s
+ N_VDD_XI13.XI24.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI13.XI27.MM25 N_XI13.XI27.CLKB_XI13.XI27.MM25_d
+ N_XI13.XI27.NET35_XI13.XI27.MM25_g N_VDD_XI13.XI27.MM25_s
+ N_VDD_XI13.XI27.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI13.XI22.MM25 N_XI13.XI22.CLKB_XI13.XI22.MM25_d
+ N_XI13.XI22.NET35_XI13.XI22.MM25_g N_VDD_XI13.XI22.MM25_s
+ N_VDD_XI13.XI22.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI13.XI21.MM25 N_XI13.XI21.CLKB_XI13.XI21.MM25_d
+ N_XI13.XI21.NET35_XI13.XI21.MM25_g N_VDD_XI13.XI21.MM25_s
+ N_VDD_XI13.XI21.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI13.XI23.MM25 N_XI13.XI23.CLKB_XI13.XI23.MM25_d
+ N_XI13.XI23.NET35_XI13.XI23.MM25_g N_VDD_XI13.XI23.MM25_s
+ N_VDD_XI13.XI23.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI13.XI19.MM25 N_XI13.XI19.CLKB_XI13.XI19.MM25_d
+ N_XI13.XI19.NET35_XI13.XI19.MM25_g N_VDD_XI13.XI19.MM25_s
+ N_VDD_XI13.XI19.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI13.XI20.MM25 N_XI13.XI20.CLKB_XI13.XI20.MM25_d
+ N_XI13.XI20.NET35_XI13.XI20.MM25_g N_VDD_XI13.XI20.MM25_s
+ N_VDD_XI13.XI20.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI13.XI18.MM25 N_XI13.XI18.CLKB_XI13.XI18.MM25_d
+ N_XI13.XI18.NET35_XI13.XI18.MM25_g N_VDD_XI13.XI18.MM25_s
+ N_VDD_XI13.XI18.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI13.XI17.MM25 N_XI13.XI17.CLKB_XI13.XI17.MM25_d
+ N_XI13.XI17.NET35_XI13.XI17.MM25_g N_VDD_XI13.XI17.MM25_s
+ N_VDD_XI13.XI17.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI13.XI0.MM25 N_XI13.XI0.CLKB_XI13.XI0.MM25_d N_XI13.XI0.NET35_XI13.XI0.MM25_g
+ N_VDD_XI13.XI0.MM25_s N_VDD_XI13.XI0.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI13.XI30.MM20 N_XI13.XI30.NET27_XI13.XI30.MM20_d N_NET382_XI13.XI30.MM20_g
+ N_VDD_XI13.XI30.MM20_s N_VDD_XI13.XI30.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI13.XI29.MM20 N_XI13.XI29.NET27_XI13.XI29.MM20_d N_NET383_XI13.XI29.MM20_g
+ N_VDD_XI13.XI29.MM20_s N_VDD_XI13.XI29.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI13.XI31.MM20 N_XI13.XI31.NET27_XI13.XI31.MM20_d N_NET384_XI13.XI31.MM20_g
+ N_VDD_XI13.XI31.MM20_s N_VDD_XI13.XI31.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI13.XI28.MM20 N_XI13.XI28.NET27_XI13.XI28.MM20_d N_NET385_XI13.XI28.MM20_g
+ N_VDD_XI13.XI28.MM20_s N_VDD_XI13.XI28.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI13.XI25.MM20 N_XI13.XI25.NET27_XI13.XI25.MM20_d N_NET386_XI13.XI25.MM20_g
+ N_VDD_XI13.XI25.MM20_s N_VDD_XI13.XI25.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI13.XI26.MM20 N_XI13.XI26.NET27_XI13.XI26.MM20_d N_NET387_XI13.XI26.MM20_g
+ N_VDD_XI13.XI26.MM20_s N_VDD_XI13.XI26.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI13.XI24.MM20 N_XI13.XI24.NET27_XI13.XI24.MM20_d N_NET388_XI13.XI24.MM20_g
+ N_VDD_XI13.XI24.MM20_s N_VDD_XI13.XI24.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI13.XI27.MM20 N_XI13.XI27.NET27_XI13.XI27.MM20_d N_NET389_XI13.XI27.MM20_g
+ N_VDD_XI13.XI27.MM20_s N_VDD_XI13.XI27.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI13.XI22.MM20 N_XI13.XI22.NET27_XI13.XI22.MM20_d N_NET390_XI13.XI22.MM20_g
+ N_VDD_XI13.XI22.MM20_s N_VDD_XI13.XI22.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI13.XI21.MM20 N_XI13.XI21.NET27_XI13.XI21.MM20_d N_NET391_XI13.XI21.MM20_g
+ N_VDD_XI13.XI21.MM20_s N_VDD_XI13.XI21.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI13.XI23.MM20 N_XI13.XI23.NET27_XI13.XI23.MM20_d N_NET392_XI13.XI23.MM20_g
+ N_VDD_XI13.XI23.MM20_s N_VDD_XI13.XI23.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI13.XI19.MM20 N_XI13.XI19.NET27_XI13.XI19.MM20_d N_NET393_XI13.XI19.MM20_g
+ N_VDD_XI13.XI19.MM20_s N_VDD_XI13.XI19.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI13.XI20.MM20 N_XI13.XI20.NET27_XI13.XI20.MM20_d N_NET394_XI13.XI20.MM20_g
+ N_VDD_XI13.XI20.MM20_s N_VDD_XI13.XI20.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI13.XI18.MM20 N_XI13.XI18.NET27_XI13.XI18.MM20_d N_NET395_XI13.XI18.MM20_g
+ N_VDD_XI13.XI18.MM20_s N_VDD_XI13.XI18.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI13.XI17.MM20 N_XI13.XI17.NET27_XI13.XI17.MM20_d N_NET396_XI13.XI17.MM20_g
+ N_VDD_XI13.XI17.MM20_s N_VDD_XI13.XI17.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI13.XI0.MM20 N_XI13.XI0.NET27_XI13.XI0.MM20_d N_NET397_XI13.XI0.MM20_g
+ N_VDD_XI13.XI0.MM20_s N_VDD_XI13.XI0.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI13.XI30.MM17 N_XI13.XI30.NET31_XI13.XI30.MM17_d
+ N_XI13.XI30.NET27_XI13.XI30.MM17_g N_VDD_XI13.XI30.MM17_s
+ N_VDD_XI13.XI30.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI13.XI29.MM17 N_XI13.XI29.NET31_XI13.XI29.MM17_d
+ N_XI13.XI29.NET27_XI13.XI29.MM17_g N_VDD_XI13.XI29.MM17_s
+ N_VDD_XI13.XI29.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI13.XI31.MM17 N_XI13.XI31.NET31_XI13.XI31.MM17_d
+ N_XI13.XI31.NET27_XI13.XI31.MM17_g N_VDD_XI13.XI31.MM17_s
+ N_VDD_XI13.XI31.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI13.XI28.MM17 N_XI13.XI28.NET31_XI13.XI28.MM17_d
+ N_XI13.XI28.NET27_XI13.XI28.MM17_g N_VDD_XI13.XI28.MM17_s
+ N_VDD_XI13.XI28.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI13.XI25.MM17 N_XI13.XI25.NET31_XI13.XI25.MM17_d
+ N_XI13.XI25.NET27_XI13.XI25.MM17_g N_VDD_XI13.XI25.MM17_s
+ N_VDD_XI13.XI25.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI13.XI26.MM17 N_XI13.XI26.NET31_XI13.XI26.MM17_d
+ N_XI13.XI26.NET27_XI13.XI26.MM17_g N_VDD_XI13.XI26.MM17_s
+ N_VDD_XI13.XI26.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI13.XI24.MM17 N_XI13.XI24.NET31_XI13.XI24.MM17_d
+ N_XI13.XI24.NET27_XI13.XI24.MM17_g N_VDD_XI13.XI24.MM17_s
+ N_VDD_XI13.XI24.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI13.XI27.MM17 N_XI13.XI27.NET31_XI13.XI27.MM17_d
+ N_XI13.XI27.NET27_XI13.XI27.MM17_g N_VDD_XI13.XI27.MM17_s
+ N_VDD_XI13.XI27.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI13.XI22.MM17 N_XI13.XI22.NET31_XI13.XI22.MM17_d
+ N_XI13.XI22.NET27_XI13.XI22.MM17_g N_VDD_XI13.XI22.MM17_s
+ N_VDD_XI13.XI22.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI13.XI21.MM17 N_XI13.XI21.NET31_XI13.XI21.MM17_d
+ N_XI13.XI21.NET27_XI13.XI21.MM17_g N_VDD_XI13.XI21.MM17_s
+ N_VDD_XI13.XI21.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI13.XI23.MM17 N_XI13.XI23.NET31_XI13.XI23.MM17_d
+ N_XI13.XI23.NET27_XI13.XI23.MM17_g N_VDD_XI13.XI23.MM17_s
+ N_VDD_XI13.XI23.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI13.XI19.MM17 N_XI13.XI19.NET31_XI13.XI19.MM17_d
+ N_XI13.XI19.NET27_XI13.XI19.MM17_g N_VDD_XI13.XI19.MM17_s
+ N_VDD_XI13.XI19.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI13.XI20.MM17 N_XI13.XI20.NET31_XI13.XI20.MM17_d
+ N_XI13.XI20.NET27_XI13.XI20.MM17_g N_VDD_XI13.XI20.MM17_s
+ N_VDD_XI13.XI20.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI13.XI18.MM17 N_XI13.XI18.NET31_XI13.XI18.MM17_d
+ N_XI13.XI18.NET27_XI13.XI18.MM17_g N_VDD_XI13.XI18.MM17_s
+ N_VDD_XI13.XI18.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI13.XI17.MM17 N_XI13.XI17.NET31_XI13.XI17.MM17_d
+ N_XI13.XI17.NET27_XI13.XI17.MM17_g N_VDD_XI13.XI17.MM17_s
+ N_VDD_XI13.XI17.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI13.XI0.MM17 N_XI13.XI0.NET31_XI13.XI0.MM17_d N_XI13.XI0.NET27_XI13.XI0.MM17_g
+ N_VDD_XI13.XI0.MM17_s N_VDD_XI13.XI0.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI13.XI30.MM27 N_XI13.XI30.NET31_XI13.XI30.MM27_d
+ N_XI13.XI30.NET35_XI13.XI30.MM27_g N_XI13.XI30.NET58_XI13.XI30.MM27_s
+ N_VDD_XI13.XI30.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=1.125e-12 AS=9.375e-13
+ PD=3e-06 PS=2.75e-06
mXI13.XI29.MM27 N_XI13.XI29.NET31_XI13.XI29.MM27_d
+ N_XI13.XI29.NET35_XI13.XI29.MM27_g N_XI13.XI29.NET58_XI13.XI29.MM27_s
+ N_VDD_XI13.XI29.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=1.125e-12 AS=9.375e-13
+ PD=3e-06 PS=2.75e-06
mXI13.XI31.MM27 N_XI13.XI31.NET31_XI13.XI31.MM27_d
+ N_XI13.XI31.NET35_XI13.XI31.MM27_g N_XI13.XI31.NET58_XI13.XI31.MM27_s
+ N_VDD_XI13.XI31.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=1.125e-12 AS=9.375e-13
+ PD=3e-06 PS=2.75e-06
mXI13.XI28.MM27 N_XI13.XI28.NET31_XI13.XI28.MM27_d
+ N_XI13.XI28.NET35_XI13.XI28.MM27_g N_XI13.XI28.NET58_XI13.XI28.MM27_s
+ N_VDD_XI13.XI28.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=1.125e-12 AS=9.375e-13
+ PD=3e-06 PS=2.75e-06
mXI13.XI25.MM27 N_XI13.XI25.NET31_XI13.XI25.MM27_d
+ N_XI13.XI25.NET35_XI13.XI25.MM27_g N_XI13.XI25.NET58_XI13.XI25.MM27_s
+ N_VDD_XI13.XI25.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=1.125e-12 AS=9.375e-13
+ PD=3e-06 PS=2.75e-06
mXI13.XI26.MM27 N_XI13.XI26.NET31_XI13.XI26.MM27_d
+ N_XI13.XI26.NET35_XI13.XI26.MM27_g N_XI13.XI26.NET58_XI13.XI26.MM27_s
+ N_VDD_XI13.XI26.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=1.125e-12 AS=9.375e-13
+ PD=3e-06 PS=2.75e-06
mXI13.XI24.MM27 N_XI13.XI24.NET31_XI13.XI24.MM27_d
+ N_XI13.XI24.NET35_XI13.XI24.MM27_g N_XI13.XI24.NET58_XI13.XI24.MM27_s
+ N_VDD_XI13.XI24.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=1.125e-12 AS=9.375e-13
+ PD=3e-06 PS=2.75e-06
mXI13.XI27.MM27 N_XI13.XI27.NET31_XI13.XI27.MM27_d
+ N_XI13.XI27.NET35_XI13.XI27.MM27_g N_XI13.XI27.NET58_XI13.XI27.MM27_s
+ N_VDD_XI13.XI27.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=1.125e-12 AS=9.375e-13
+ PD=3e-06 PS=2.75e-06
mXI13.XI22.MM27 N_XI13.XI22.NET31_XI13.XI22.MM27_d
+ N_XI13.XI22.NET35_XI13.XI22.MM27_g N_XI13.XI22.NET58_XI13.XI22.MM27_s
+ N_VDD_XI13.XI22.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=1.125e-12 AS=9.375e-13
+ PD=3e-06 PS=2.75e-06
mXI13.XI21.MM27 N_XI13.XI21.NET31_XI13.XI21.MM27_d
+ N_XI13.XI21.NET35_XI13.XI21.MM27_g N_XI13.XI21.NET58_XI13.XI21.MM27_s
+ N_VDD_XI13.XI21.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=1.125e-12 AS=9.375e-13
+ PD=3e-06 PS=2.75e-06
mXI13.XI23.MM27 N_XI13.XI23.NET31_XI13.XI23.MM27_d
+ N_XI13.XI23.NET35_XI13.XI23.MM27_g N_XI13.XI23.NET58_XI13.XI23.MM27_s
+ N_VDD_XI13.XI23.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=1.125e-12 AS=9.375e-13
+ PD=3e-06 PS=2.75e-06
mXI13.XI19.MM27 N_XI13.XI19.NET31_XI13.XI19.MM27_d
+ N_XI13.XI19.NET35_XI13.XI19.MM27_g N_XI13.XI19.NET58_XI13.XI19.MM27_s
+ N_VDD_XI13.XI19.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=1.125e-12 AS=9.375e-13
+ PD=3e-06 PS=2.75e-06
mXI13.XI20.MM27 N_XI13.XI20.NET31_XI13.XI20.MM27_d
+ N_XI13.XI20.NET35_XI13.XI20.MM27_g N_XI13.XI20.NET58_XI13.XI20.MM27_s
+ N_VDD_XI13.XI20.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=1.125e-12 AS=9.375e-13
+ PD=3e-06 PS=2.75e-06
mXI13.XI18.MM27 N_XI13.XI18.NET31_XI13.XI18.MM27_d
+ N_XI13.XI18.NET35_XI13.XI18.MM27_g N_XI13.XI18.NET58_XI13.XI18.MM27_s
+ N_VDD_XI13.XI18.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=1.125e-12 AS=9.375e-13
+ PD=3e-06 PS=2.75e-06
mXI13.XI17.MM27 N_XI13.XI17.NET31_XI13.XI17.MM27_d
+ N_XI13.XI17.NET35_XI13.XI17.MM27_g N_XI13.XI17.NET58_XI13.XI17.MM27_s
+ N_VDD_XI13.XI17.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=1.125e-12 AS=9.375e-13
+ PD=3e-06 PS=2.75e-06
mXI13.XI0.MM27 N_XI13.XI0.NET31_XI13.XI0.MM27_d N_XI13.XI0.NET35_XI13.XI0.MM27_g
+ N_XI13.XI0.NET58_XI13.XI0.MM27_s N_VDD_XI13.XI0.XI0.MM1_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.125e-12 AS=9.375e-13 PD=3e-06 PS=2.75e-06
mXI13.XI30.MM3 N_XI13.XI30.NET15_XI13.XI30.MM3_d
+ N_XI13.XI30.NET58_XI13.XI30.MM3_g N_VDD_XI13.XI30.MM3_s
+ N_VDD_XI13.XI30.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI13.XI29.MM3 N_XI13.XI29.NET15_XI13.XI29.MM3_d
+ N_XI13.XI29.NET58_XI13.XI29.MM3_g N_VDD_XI13.XI29.MM3_s
+ N_VDD_XI13.XI29.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI13.XI31.MM3 N_XI13.XI31.NET15_XI13.XI31.MM3_d
+ N_XI13.XI31.NET58_XI13.XI31.MM3_g N_VDD_XI13.XI31.MM3_s
+ N_VDD_XI13.XI31.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI13.XI28.MM3 N_XI13.XI28.NET15_XI13.XI28.MM3_d
+ N_XI13.XI28.NET58_XI13.XI28.MM3_g N_VDD_XI13.XI28.MM3_s
+ N_VDD_XI13.XI28.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI13.XI25.MM3 N_XI13.XI25.NET15_XI13.XI25.MM3_d
+ N_XI13.XI25.NET58_XI13.XI25.MM3_g N_VDD_XI13.XI25.MM3_s
+ N_VDD_XI13.XI25.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI13.XI26.MM3 N_XI13.XI26.NET15_XI13.XI26.MM3_d
+ N_XI13.XI26.NET58_XI13.XI26.MM3_g N_VDD_XI13.XI26.MM3_s
+ N_VDD_XI13.XI26.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI13.XI24.MM3 N_XI13.XI24.NET15_XI13.XI24.MM3_d
+ N_XI13.XI24.NET58_XI13.XI24.MM3_g N_VDD_XI13.XI24.MM3_s
+ N_VDD_XI13.XI24.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI13.XI27.MM3 N_XI13.XI27.NET15_XI13.XI27.MM3_d
+ N_XI13.XI27.NET58_XI13.XI27.MM3_g N_VDD_XI13.XI27.MM3_s
+ N_VDD_XI13.XI27.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI13.XI22.MM3 N_XI13.XI22.NET15_XI13.XI22.MM3_d
+ N_XI13.XI22.NET58_XI13.XI22.MM3_g N_VDD_XI13.XI22.MM3_s
+ N_VDD_XI13.XI22.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI13.XI21.MM3 N_XI13.XI21.NET15_XI13.XI21.MM3_d
+ N_XI13.XI21.NET58_XI13.XI21.MM3_g N_VDD_XI13.XI21.MM3_s
+ N_VDD_XI13.XI21.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI13.XI23.MM3 N_XI13.XI23.NET15_XI13.XI23.MM3_d
+ N_XI13.XI23.NET58_XI13.XI23.MM3_g N_VDD_XI13.XI23.MM3_s
+ N_VDD_XI13.XI23.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI13.XI19.MM3 N_XI13.XI19.NET15_XI13.XI19.MM3_d
+ N_XI13.XI19.NET58_XI13.XI19.MM3_g N_VDD_XI13.XI19.MM3_s
+ N_VDD_XI13.XI19.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI13.XI20.MM3 N_XI13.XI20.NET15_XI13.XI20.MM3_d
+ N_XI13.XI20.NET58_XI13.XI20.MM3_g N_VDD_XI13.XI20.MM3_s
+ N_VDD_XI13.XI20.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI13.XI18.MM3 N_XI13.XI18.NET15_XI13.XI18.MM3_d
+ N_XI13.XI18.NET58_XI13.XI18.MM3_g N_VDD_XI13.XI18.MM3_s
+ N_VDD_XI13.XI18.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI13.XI17.MM3 N_XI13.XI17.NET15_XI13.XI17.MM3_d
+ N_XI13.XI17.NET58_XI13.XI17.MM3_g N_VDD_XI13.XI17.MM3_s
+ N_VDD_XI13.XI17.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI13.XI0.MM3 N_XI13.XI0.NET15_XI13.XI0.MM3_d N_XI13.XI0.NET58_XI13.XI0.MM3_g
+ N_VDD_XI13.XI0.MM3_s N_VDD_XI13.XI0.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI13.XI30.MM1 N_XI13.XI30.NET54_XI13.XI30.MM1_d
+ N_XI13.XI30.NET15_XI13.XI30.MM1_g N_VDD_XI13.XI30.MM1_s
+ N_VDD_XI13.XI30.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI13.XI29.MM1 N_XI13.XI29.NET54_XI13.XI29.MM1_d
+ N_XI13.XI29.NET15_XI13.XI29.MM1_g N_VDD_XI13.XI29.MM1_s
+ N_VDD_XI13.XI29.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI13.XI31.MM1 N_XI13.XI31.NET54_XI13.XI31.MM1_d
+ N_XI13.XI31.NET15_XI13.XI31.MM1_g N_VDD_XI13.XI31.MM1_s
+ N_VDD_XI13.XI31.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI13.XI28.MM1 N_XI13.XI28.NET54_XI13.XI28.MM1_d
+ N_XI13.XI28.NET15_XI13.XI28.MM1_g N_VDD_XI13.XI28.MM1_s
+ N_VDD_XI13.XI28.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI13.XI25.MM1 N_XI13.XI25.NET54_XI13.XI25.MM1_d
+ N_XI13.XI25.NET15_XI13.XI25.MM1_g N_VDD_XI13.XI25.MM1_s
+ N_VDD_XI13.XI25.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI13.XI26.MM1 N_XI13.XI26.NET54_XI13.XI26.MM1_d
+ N_XI13.XI26.NET15_XI13.XI26.MM1_g N_VDD_XI13.XI26.MM1_s
+ N_VDD_XI13.XI26.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI13.XI24.MM1 N_XI13.XI24.NET54_XI13.XI24.MM1_d
+ N_XI13.XI24.NET15_XI13.XI24.MM1_g N_VDD_XI13.XI24.MM1_s
+ N_VDD_XI13.XI24.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI13.XI27.MM1 N_XI13.XI27.NET54_XI13.XI27.MM1_d
+ N_XI13.XI27.NET15_XI13.XI27.MM1_g N_VDD_XI13.XI27.MM1_s
+ N_VDD_XI13.XI27.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI13.XI22.MM1 N_XI13.XI22.NET54_XI13.XI22.MM1_d
+ N_XI13.XI22.NET15_XI13.XI22.MM1_g N_VDD_XI13.XI22.MM1_s
+ N_VDD_XI13.XI22.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI13.XI21.MM1 N_XI13.XI21.NET54_XI13.XI21.MM1_d
+ N_XI13.XI21.NET15_XI13.XI21.MM1_g N_VDD_XI13.XI21.MM1_s
+ N_VDD_XI13.XI21.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI13.XI23.MM1 N_XI13.XI23.NET54_XI13.XI23.MM1_d
+ N_XI13.XI23.NET15_XI13.XI23.MM1_g N_VDD_XI13.XI23.MM1_s
+ N_VDD_XI13.XI23.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI13.XI19.MM1 N_XI13.XI19.NET54_XI13.XI19.MM1_d
+ N_XI13.XI19.NET15_XI13.XI19.MM1_g N_VDD_XI13.XI19.MM1_s
+ N_VDD_XI13.XI19.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI13.XI20.MM1 N_XI13.XI20.NET54_XI13.XI20.MM1_d
+ N_XI13.XI20.NET15_XI13.XI20.MM1_g N_VDD_XI13.XI20.MM1_s
+ N_VDD_XI13.XI20.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI13.XI18.MM1 N_XI13.XI18.NET54_XI13.XI18.MM1_d
+ N_XI13.XI18.NET15_XI13.XI18.MM1_g N_VDD_XI13.XI18.MM1_s
+ N_VDD_XI13.XI18.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI13.XI17.MM1 N_XI13.XI17.NET54_XI13.XI17.MM1_d
+ N_XI13.XI17.NET15_XI13.XI17.MM1_g N_VDD_XI13.XI17.MM1_s
+ N_VDD_XI13.XI17.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI13.XI0.MM1 N_XI13.XI0.NET54_XI13.XI0.MM1_d N_XI13.XI0.NET15_XI13.XI0.MM1_g
+ N_VDD_XI13.XI0.MM1_s N_VDD_XI13.XI0.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI13.XI30.MM35 N_XI13.XI30.NET58_XI13.XI30.MM35_d
+ N_XI13.XI30.CLKB_XI13.XI30.MM35_g N_XI13.XI30.NET54_XI13.XI30.MM35_s
+ N_VDD_XI13.XI30.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI13.XI29.MM35 N_XI13.XI29.NET58_XI13.XI29.MM35_d
+ N_XI13.XI29.CLKB_XI13.XI29.MM35_g N_XI13.XI29.NET54_XI13.XI29.MM35_s
+ N_VDD_XI13.XI29.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI13.XI31.MM35 N_XI13.XI31.NET58_XI13.XI31.MM35_d
+ N_XI13.XI31.CLKB_XI13.XI31.MM35_g N_XI13.XI31.NET54_XI13.XI31.MM35_s
+ N_VDD_XI13.XI31.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI13.XI28.MM35 N_XI13.XI28.NET58_XI13.XI28.MM35_d
+ N_XI13.XI28.CLKB_XI13.XI28.MM35_g N_XI13.XI28.NET54_XI13.XI28.MM35_s
+ N_VDD_XI13.XI28.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI13.XI25.MM35 N_XI13.XI25.NET58_XI13.XI25.MM35_d
+ N_XI13.XI25.CLKB_XI13.XI25.MM35_g N_XI13.XI25.NET54_XI13.XI25.MM35_s
+ N_VDD_XI13.XI25.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI13.XI26.MM35 N_XI13.XI26.NET58_XI13.XI26.MM35_d
+ N_XI13.XI26.CLKB_XI13.XI26.MM35_g N_XI13.XI26.NET54_XI13.XI26.MM35_s
+ N_VDD_XI13.XI26.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI13.XI24.MM35 N_XI13.XI24.NET58_XI13.XI24.MM35_d
+ N_XI13.XI24.CLKB_XI13.XI24.MM35_g N_XI13.XI24.NET54_XI13.XI24.MM35_s
+ N_VDD_XI13.XI24.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI13.XI27.MM35 N_XI13.XI27.NET58_XI13.XI27.MM35_d
+ N_XI13.XI27.CLKB_XI13.XI27.MM35_g N_XI13.XI27.NET54_XI13.XI27.MM35_s
+ N_VDD_XI13.XI27.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI13.XI22.MM35 N_XI13.XI22.NET58_XI13.XI22.MM35_d
+ N_XI13.XI22.CLKB_XI13.XI22.MM35_g N_XI13.XI22.NET54_XI13.XI22.MM35_s
+ N_VDD_XI13.XI22.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI13.XI21.MM35 N_XI13.XI21.NET58_XI13.XI21.MM35_d
+ N_XI13.XI21.CLKB_XI13.XI21.MM35_g N_XI13.XI21.NET54_XI13.XI21.MM35_s
+ N_VDD_XI13.XI21.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI13.XI23.MM35 N_XI13.XI23.NET58_XI13.XI23.MM35_d
+ N_XI13.XI23.CLKB_XI13.XI23.MM35_g N_XI13.XI23.NET54_XI13.XI23.MM35_s
+ N_VDD_XI13.XI23.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI13.XI19.MM35 N_XI13.XI19.NET58_XI13.XI19.MM35_d
+ N_XI13.XI19.CLKB_XI13.XI19.MM35_g N_XI13.XI19.NET54_XI13.XI19.MM35_s
+ N_VDD_XI13.XI19.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI13.XI20.MM35 N_XI13.XI20.NET58_XI13.XI20.MM35_d
+ N_XI13.XI20.CLKB_XI13.XI20.MM35_g N_XI13.XI20.NET54_XI13.XI20.MM35_s
+ N_VDD_XI13.XI20.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI13.XI18.MM35 N_XI13.XI18.NET58_XI13.XI18.MM35_d
+ N_XI13.XI18.CLKB_XI13.XI18.MM35_g N_XI13.XI18.NET54_XI13.XI18.MM35_s
+ N_VDD_XI13.XI18.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI13.XI17.MM35 N_XI13.XI17.NET58_XI13.XI17.MM35_d
+ N_XI13.XI17.CLKB_XI13.XI17.MM35_g N_XI13.XI17.NET54_XI13.XI17.MM35_s
+ N_VDD_XI13.XI17.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI13.XI0.MM35 N_XI13.XI0.NET58_XI13.XI0.MM35_d N_XI13.XI0.CLKB_XI13.XI0.MM35_g
+ N_XI13.XI0.NET54_XI13.XI0.MM35_s N_VDD_XI13.XI0.XI0.MM1_b P_18 L=1.8e-07
+ W=1.5e-06 AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI13.XI30.MM37 N_XI13.XI30.NET15_XI13.XI30.MM37_d
+ N_XI13.XI30.CLKB_XI13.XI30.MM37_g N_XI13.XI30.NET14_XI13.XI30.MM37_s
+ N_VDD_XI13.XI30.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=1.125e-12 AS=9.375e-13
+ PD=3e-06 PS=2.75e-06
mXI13.XI29.MM37 N_XI13.XI29.NET15_XI13.XI29.MM37_d
+ N_XI13.XI29.CLKB_XI13.XI29.MM37_g N_XI13.XI29.NET14_XI13.XI29.MM37_s
+ N_VDD_XI13.XI29.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=1.125e-12 AS=9.375e-13
+ PD=3e-06 PS=2.75e-06
mXI13.XI31.MM37 N_XI13.XI31.NET15_XI13.XI31.MM37_d
+ N_XI13.XI31.CLKB_XI13.XI31.MM37_g N_XI13.XI31.NET14_XI13.XI31.MM37_s
+ N_VDD_XI13.XI31.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=1.125e-12 AS=9.375e-13
+ PD=3e-06 PS=2.75e-06
mXI13.XI28.MM37 N_XI13.XI28.NET15_XI13.XI28.MM37_d
+ N_XI13.XI28.CLKB_XI13.XI28.MM37_g N_XI13.XI28.NET14_XI13.XI28.MM37_s
+ N_VDD_XI13.XI28.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=1.125e-12 AS=9.375e-13
+ PD=3e-06 PS=2.75e-06
mXI13.XI25.MM37 N_XI13.XI25.NET15_XI13.XI25.MM37_d
+ N_XI13.XI25.CLKB_XI13.XI25.MM37_g N_XI13.XI25.NET14_XI13.XI25.MM37_s
+ N_VDD_XI13.XI25.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=1.125e-12 AS=9.375e-13
+ PD=3e-06 PS=2.75e-06
mXI13.XI26.MM37 N_XI13.XI26.NET15_XI13.XI26.MM37_d
+ N_XI13.XI26.CLKB_XI13.XI26.MM37_g N_XI13.XI26.NET14_XI13.XI26.MM37_s
+ N_VDD_XI13.XI26.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=1.125e-12 AS=9.375e-13
+ PD=3e-06 PS=2.75e-06
mXI13.XI24.MM37 N_XI13.XI24.NET15_XI13.XI24.MM37_d
+ N_XI13.XI24.CLKB_XI13.XI24.MM37_g N_XI13.XI24.NET14_XI13.XI24.MM37_s
+ N_VDD_XI13.XI24.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=1.125e-12 AS=9.375e-13
+ PD=3e-06 PS=2.75e-06
mXI13.XI27.MM37 N_XI13.XI27.NET15_XI13.XI27.MM37_d
+ N_XI13.XI27.CLKB_XI13.XI27.MM37_g N_XI13.XI27.NET14_XI13.XI27.MM37_s
+ N_VDD_XI13.XI27.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=1.125e-12 AS=9.375e-13
+ PD=3e-06 PS=2.75e-06
mXI13.XI22.MM37 N_XI13.XI22.NET15_XI13.XI22.MM37_d
+ N_XI13.XI22.CLKB_XI13.XI22.MM37_g N_XI13.XI22.NET14_XI13.XI22.MM37_s
+ N_VDD_XI13.XI22.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=1.125e-12 AS=9.375e-13
+ PD=3e-06 PS=2.75e-06
mXI13.XI21.MM37 N_XI13.XI21.NET15_XI13.XI21.MM37_d
+ N_XI13.XI21.CLKB_XI13.XI21.MM37_g N_XI13.XI21.NET14_XI13.XI21.MM37_s
+ N_VDD_XI13.XI21.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=1.125e-12 AS=9.375e-13
+ PD=3e-06 PS=2.75e-06
mXI13.XI23.MM37 N_XI13.XI23.NET15_XI13.XI23.MM37_d
+ N_XI13.XI23.CLKB_XI13.XI23.MM37_g N_XI13.XI23.NET14_XI13.XI23.MM37_s
+ N_VDD_XI13.XI23.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=1.125e-12 AS=9.375e-13
+ PD=3e-06 PS=2.75e-06
mXI13.XI19.MM37 N_XI13.XI19.NET15_XI13.XI19.MM37_d
+ N_XI13.XI19.CLKB_XI13.XI19.MM37_g N_XI13.XI19.NET14_XI13.XI19.MM37_s
+ N_VDD_XI13.XI19.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=1.125e-12 AS=9.375e-13
+ PD=3e-06 PS=2.75e-06
mXI13.XI20.MM37 N_XI13.XI20.NET15_XI13.XI20.MM37_d
+ N_XI13.XI20.CLKB_XI13.XI20.MM37_g N_XI13.XI20.NET14_XI13.XI20.MM37_s
+ N_VDD_XI13.XI20.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=1.125e-12 AS=9.375e-13
+ PD=3e-06 PS=2.75e-06
mXI13.XI18.MM37 N_XI13.XI18.NET15_XI13.XI18.MM37_d
+ N_XI13.XI18.CLKB_XI13.XI18.MM37_g N_XI13.XI18.NET14_XI13.XI18.MM37_s
+ N_VDD_XI13.XI18.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=1.125e-12 AS=9.375e-13
+ PD=3e-06 PS=2.75e-06
mXI13.XI17.MM37 N_XI13.XI17.NET15_XI13.XI17.MM37_d
+ N_XI13.XI17.CLKB_XI13.XI17.MM37_g N_XI13.XI17.NET14_XI13.XI17.MM37_s
+ N_VDD_XI13.XI17.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=1.125e-12 AS=9.375e-13
+ PD=3e-06 PS=2.75e-06
mXI13.XI0.MM37 N_XI13.XI0.NET15_XI13.XI0.MM37_d N_XI13.XI0.CLKB_XI13.XI0.MM37_g
+ N_XI13.XI0.NET14_XI13.XI0.MM37_s N_VDD_XI13.XI0.XI0.MM1_b P_18 L=1.8e-07
+ W=1.5e-06 AD=1.125e-12 AS=9.375e-13 PD=3e-06 PS=2.75e-06
mXI13.XI30.MM13 N_MAX15_XI13.XI30.MM13_d N_XI13.XI30.NET14_XI13.XI30.MM13_g
+ N_VDD_XI13.XI30.MM13_s N_VDD_XI13.XI30.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI13.XI29.MM13 N_MAX14_XI13.XI29.MM13_d N_XI13.XI29.NET14_XI13.XI29.MM13_g
+ N_VDD_XI13.XI29.MM13_s N_VDD_XI13.XI29.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI13.XI31.MM13 N_MAX13_XI13.XI31.MM13_d N_XI13.XI31.NET14_XI13.XI31.MM13_g
+ N_VDD_XI13.XI31.MM13_s N_VDD_XI13.XI31.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI13.XI28.MM13 N_MAX12_XI13.XI28.MM13_d N_XI13.XI28.NET14_XI13.XI28.MM13_g
+ N_VDD_XI13.XI28.MM13_s N_VDD_XI13.XI28.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI13.XI25.MM13 N_MAX11_XI13.XI25.MM13_d N_XI13.XI25.NET14_XI13.XI25.MM13_g
+ N_VDD_XI13.XI25.MM13_s N_VDD_XI13.XI25.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI13.XI26.MM13 N_MAX10_XI13.XI26.MM13_d N_XI13.XI26.NET14_XI13.XI26.MM13_g
+ N_VDD_XI13.XI26.MM13_s N_VDD_XI13.XI26.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI13.XI24.MM13 N_MAX9_XI13.XI24.MM13_d N_XI13.XI24.NET14_XI13.XI24.MM13_g
+ N_VDD_XI13.XI24.MM13_s N_VDD_XI13.XI24.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI13.XI27.MM13 N_MAX8_XI13.XI27.MM13_d N_XI13.XI27.NET14_XI13.XI27.MM13_g
+ N_VDD_XI13.XI27.MM13_s N_VDD_XI13.XI27.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI13.XI22.MM13 N_MAX7_XI13.XI22.MM13_d N_XI13.XI22.NET14_XI13.XI22.MM13_g
+ N_VDD_XI13.XI22.MM13_s N_VDD_XI13.XI22.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI13.XI21.MM13 N_MAX6_XI13.XI21.MM13_d N_XI13.XI21.NET14_XI13.XI21.MM13_g
+ N_VDD_XI13.XI21.MM13_s N_VDD_XI13.XI21.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI13.XI23.MM13 N_MAX5_XI13.XI23.MM13_d N_XI13.XI23.NET14_XI13.XI23.MM13_g
+ N_VDD_XI13.XI23.MM13_s N_VDD_XI13.XI23.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI13.XI19.MM13 N_MAX4_XI13.XI19.MM13_d N_XI13.XI19.NET14_XI13.XI19.MM13_g
+ N_VDD_XI13.XI19.MM13_s N_VDD_XI13.XI19.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI13.XI20.MM13 N_MAX3_XI13.XI20.MM13_d N_XI13.XI20.NET14_XI13.XI20.MM13_g
+ N_VDD_XI13.XI20.MM13_s N_VDD_XI13.XI20.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI13.XI18.MM13 N_MAX2_XI13.XI18.MM13_d N_XI13.XI18.NET14_XI13.XI18.MM13_g
+ N_VDD_XI13.XI18.MM13_s N_VDD_XI13.XI18.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI13.XI17.MM13 N_MAX1_XI13.XI17.MM13_d N_XI13.XI17.NET14_XI13.XI17.MM13_g
+ N_VDD_XI13.XI17.MM13_s N_VDD_XI13.XI17.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI13.XI0.MM13 N_MAX0_XI13.XI0.MM13_d N_XI13.XI0.NET14_XI13.XI0.MM13_g
+ N_VDD_XI13.XI0.MM13_s N_VDD_XI13.XI0.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI13.XI30.MM14 N_XI13.BAR_Q16_XI13.XI30.MM14_d N_MAX15_XI13.XI30.MM14_g
+ N_VDD_XI13.XI30.MM14_s N_VDD_XI13.XI30.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI13.XI29.MM14 N_XI13.BAR_Q15_XI13.XI29.MM14_d N_MAX14_XI13.XI29.MM14_g
+ N_VDD_XI13.XI29.MM14_s N_VDD_XI13.XI29.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI13.XI31.MM14 N_XI13.BAR_Q14_XI13.XI31.MM14_d N_MAX13_XI13.XI31.MM14_g
+ N_VDD_XI13.XI31.MM14_s N_VDD_XI13.XI31.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI13.XI28.MM14 N_XI13.BAR_Q13_XI13.XI28.MM14_d N_MAX12_XI13.XI28.MM14_g
+ N_VDD_XI13.XI28.MM14_s N_VDD_XI13.XI28.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI13.XI25.MM14 N_XI13.BAR_Q12_XI13.XI25.MM14_d N_MAX11_XI13.XI25.MM14_g
+ N_VDD_XI13.XI25.MM14_s N_VDD_XI13.XI25.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI13.XI26.MM14 N_XI13.BAR_Q11_XI13.XI26.MM14_d N_MAX10_XI13.XI26.MM14_g
+ N_VDD_XI13.XI26.MM14_s N_VDD_XI13.XI26.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI13.XI24.MM14 N_XI13.BAR_Q10_XI13.XI24.MM14_d N_MAX9_XI13.XI24.MM14_g
+ N_VDD_XI13.XI24.MM14_s N_VDD_XI13.XI24.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI13.XI27.MM14 N_XI13.BAR_Q9_XI13.XI27.MM14_d N_MAX8_XI13.XI27.MM14_g
+ N_VDD_XI13.XI27.MM14_s N_VDD_XI13.XI27.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI13.XI22.MM14 N_XI13.BAR_Q8_XI13.XI22.MM14_d N_MAX7_XI13.XI22.MM14_g
+ N_VDD_XI13.XI22.MM14_s N_VDD_XI13.XI22.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI13.XI21.MM14 N_XI13.BAR_Q7_XI13.XI21.MM14_d N_MAX6_XI13.XI21.MM14_g
+ N_VDD_XI13.XI21.MM14_s N_VDD_XI13.XI21.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI13.XI23.MM14 N_XI13.BAR_Q6_XI13.XI23.MM14_d N_MAX5_XI13.XI23.MM14_g
+ N_VDD_XI13.XI23.MM14_s N_VDD_XI13.XI23.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI13.XI19.MM14 N_XI13.BAR_Q5_XI13.XI19.MM14_d N_MAX4_XI13.XI19.MM14_g
+ N_VDD_XI13.XI19.MM14_s N_VDD_XI13.XI19.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI13.XI20.MM14 N_XI13.BAR_Q4_XI13.XI20.MM14_d N_MAX3_XI13.XI20.MM14_g
+ N_VDD_XI13.XI20.MM14_s N_VDD_XI13.XI20.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI13.XI18.MM14 N_XI13.BAR_Q3_XI13.XI18.MM14_d N_MAX2_XI13.XI18.MM14_g
+ N_VDD_XI13.XI18.MM14_s N_VDD_XI13.XI18.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI13.XI17.MM14 N_XI13.BAR_Q2_XI13.XI17.MM14_d N_MAX1_XI13.XI17.MM14_g
+ N_VDD_XI13.XI17.MM14_s N_VDD_XI13.XI17.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI13.XI0.MM14 N_XI13.BAR_Q1_XI13.XI0.MM14_d N_MAX0_XI13.XI0.MM14_g
+ N_VDD_XI13.XI0.MM14_s N_VDD_XI13.XI0.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06
+ AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
mXI13.XI30.MM39 N_XI13.XI30.NET14_XI13.XI30.MM39_d
+ N_XI13.XI30.NET35_XI13.XI30.MM39_g N_XI13.BAR_Q16_XI13.XI30.MM39_s
+ N_VDD_XI13.XI30.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI13.XI29.MM39 N_XI13.XI29.NET14_XI13.XI29.MM39_d
+ N_XI13.XI29.NET35_XI13.XI29.MM39_g N_XI13.BAR_Q15_XI13.XI29.MM39_s
+ N_VDD_XI13.XI29.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI13.XI31.MM39 N_XI13.XI31.NET14_XI13.XI31.MM39_d
+ N_XI13.XI31.NET35_XI13.XI31.MM39_g N_XI13.BAR_Q14_XI13.XI31.MM39_s
+ N_VDD_XI13.XI31.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI13.XI28.MM39 N_XI13.XI28.NET14_XI13.XI28.MM39_d
+ N_XI13.XI28.NET35_XI13.XI28.MM39_g N_XI13.BAR_Q13_XI13.XI28.MM39_s
+ N_VDD_XI13.XI28.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI13.XI25.MM39 N_XI13.XI25.NET14_XI13.XI25.MM39_d
+ N_XI13.XI25.NET35_XI13.XI25.MM39_g N_XI13.BAR_Q12_XI13.XI25.MM39_s
+ N_VDD_XI13.XI25.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI13.XI26.MM39 N_XI13.XI26.NET14_XI13.XI26.MM39_d
+ N_XI13.XI26.NET35_XI13.XI26.MM39_g N_XI13.BAR_Q11_XI13.XI26.MM39_s
+ N_VDD_XI13.XI26.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI13.XI24.MM39 N_XI13.XI24.NET14_XI13.XI24.MM39_d
+ N_XI13.XI24.NET35_XI13.XI24.MM39_g N_XI13.BAR_Q10_XI13.XI24.MM39_s
+ N_VDD_XI13.XI24.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI13.XI27.MM39 N_XI13.XI27.NET14_XI13.XI27.MM39_d
+ N_XI13.XI27.NET35_XI13.XI27.MM39_g N_XI13.BAR_Q9_XI13.XI27.MM39_s
+ N_VDD_XI13.XI27.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI13.XI22.MM39 N_XI13.XI22.NET14_XI13.XI22.MM39_d
+ N_XI13.XI22.NET35_XI13.XI22.MM39_g N_XI13.BAR_Q8_XI13.XI22.MM39_s
+ N_VDD_XI13.XI22.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI13.XI21.MM39 N_XI13.XI21.NET14_XI13.XI21.MM39_d
+ N_XI13.XI21.NET35_XI13.XI21.MM39_g N_XI13.BAR_Q7_XI13.XI21.MM39_s
+ N_VDD_XI13.XI21.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI13.XI23.MM39 N_XI13.XI23.NET14_XI13.XI23.MM39_d
+ N_XI13.XI23.NET35_XI13.XI23.MM39_g N_XI13.BAR_Q6_XI13.XI23.MM39_s
+ N_VDD_XI13.XI23.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI13.XI19.MM39 N_XI13.XI19.NET14_XI13.XI19.MM39_d
+ N_XI13.XI19.NET35_XI13.XI19.MM39_g N_XI13.BAR_Q5_XI13.XI19.MM39_s
+ N_VDD_XI13.XI19.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI13.XI20.MM39 N_XI13.XI20.NET14_XI13.XI20.MM39_d
+ N_XI13.XI20.NET35_XI13.XI20.MM39_g N_XI13.BAR_Q4_XI13.XI20.MM39_s
+ N_VDD_XI13.XI20.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI13.XI18.MM39 N_XI13.XI18.NET14_XI13.XI18.MM39_d
+ N_XI13.XI18.NET35_XI13.XI18.MM39_g N_XI13.BAR_Q3_XI13.XI18.MM39_s
+ N_VDD_XI13.XI18.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI13.XI17.MM39 N_XI13.XI17.NET14_XI13.XI17.MM39_d
+ N_XI13.XI17.NET35_XI13.XI17.MM39_g N_XI13.BAR_Q2_XI13.XI17.MM39_s
+ N_VDD_XI13.XI17.XI0.MM1_b P_18 L=1.8e-07 W=1.5e-06 AD=9.375e-13 AS=1.125e-12
+ PD=2.75e-06 PS=3e-06
mXI13.XI0.MM39 N_XI13.XI0.NET14_XI13.XI0.MM39_d N_XI13.XI0.NET35_XI13.XI0.MM39_g
+ N_XI13.BAR_Q1_XI13.XI0.MM39_s N_VDD_XI13.XI0.XI0.MM1_b P_18 L=1.8e-07
+ W=1.5e-06 AD=9.375e-13 AS=1.125e-12 PD=2.75e-06 PS=3e-06
*
.include "acc_min_max.pex.sp.ACC_MIN_MAX.pxi"
*
.ends
*
*
